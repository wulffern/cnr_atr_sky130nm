magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1152 2025
<< ndiff >>
rect 416 45 608 117
rect 416 117 608 981
rect 416 981 608 1053
rect 416 1053 608 1917
rect 416 1917 608 1989
<< ptap >>
rect -96 -36 96 45
rect 1056 -36 1248 45
rect -96 45 96 117
rect 1056 45 1248 117
rect -96 117 96 981
rect 1056 117 1248 981
rect -96 981 96 1053
rect 1056 981 1248 1053
rect -96 1053 96 1917
rect 1056 1053 1248 1917
rect -96 1917 96 1989
rect 1056 1917 1248 1989
rect -96 1989 96 2070
rect 1056 1989 1248 2070
<< poly >>
rect 352 -18 864 27
rect 352 135 864 963
rect 352 1071 864 1899
rect 352 2007 864 2052
rect 800 117 864 981
rect 800 981 864 1053
rect 800 1053 864 1917
<< locali >>
rect 800 1053 864 1917
rect -96 -36 96 45
rect 1056 -36 1248 45
rect -96 45 96 117
rect 288 45 608 117
rect 288 45 608 117
rect 1056 45 1248 117
rect -96 117 96 981
rect 288 117 352 981
rect 800 117 864 981
rect 1056 117 1248 981
rect -96 981 96 1053
rect 1056 981 1248 1053
rect 288 981 352 1053
rect 416 981 608 1053
rect 416 981 608 1053
rect 800 981 864 1053
rect 1056 981 1248 1053
rect -96 1053 96 1917
rect 288 1053 352 1917
rect 800 1053 864 1917
rect 1056 1053 1248 1917
rect -96 1917 96 1989
rect 288 1917 608 1989
rect 1056 1917 1248 1989
rect -96 1989 96 2070
rect 1056 1989 1248 2070
<< pcontact >>
rect 810 333 853 549
rect 810 549 853 765
rect 810 765 853 981
rect 810 981 853 999
rect 810 999 853 1017
rect 810 1017 853 1035
rect 810 1035 853 1053
rect 810 1053 853 1269
rect 810 1269 853 1485
rect 810 1485 853 1701
<< ptapc >>
rect -32 45 32 117
rect 1120 45 1184 117
rect -32 117 32 981
rect 1120 117 1184 981
rect -32 981 32 1053
rect 1120 981 1184 1053
rect -32 1053 32 1917
rect 1120 1053 1184 1917
rect -32 1917 32 1989
rect 1120 1917 1184 1989
<< ndcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 448 999 480 1017
rect 448 1017 480 1035
rect 480 999 544 1017
rect 480 1017 544 1035
rect 544 999 576 1017
rect 544 1017 576 1035
rect 448 1935 480 1953
rect 448 1953 480 1971
rect 480 1935 544 1953
rect 480 1953 544 1971
rect 544 1935 576 1953
rect 544 1953 576 1971
<< pwell >>
rect -184 -124 1336 2158
<< labels >>
flabel locali s 800 1053 864 1917 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 608 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1056 981 1248 1053 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 981 608 1053 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 2025
<< end >>
