magic
tech sky130B
magscale 1 2
timestamp 1695852000
<< checkpaint >>
rect 0 0 1728 2030
<< ndiff >>
rect 416 50 1184 122
rect 416 122 1184 986
rect 416 986 1184 1058
rect 416 1058 1184 1922
rect 416 1922 1184 1994
<< ptap >>
rect -96 -36 96 50
rect 1632 -36 1824 50
rect -96 50 96 122
rect 1632 50 1824 122
rect -96 122 96 986
rect 1632 122 1824 986
rect -96 986 96 1058
rect 1632 986 1824 1058
rect -96 1058 96 1922
rect 1632 1058 1824 1922
rect -96 1922 96 1994
rect 1632 1922 1824 1994
rect -96 1994 96 2080
rect 1632 1994 1824 2080
<< poly >>
rect 352 -18 1440 32
rect 352 140 1440 968
rect 352 1076 1440 1904
rect 352 2012 1440 2062
rect 1376 122 1440 986
rect 1376 986 1440 1058
rect 1376 1058 1440 1922
<< locali >>
rect 1376 1058 1440 1922
rect -96 -36 96 50
rect 1632 -36 1824 50
rect -96 50 96 122
rect 288 50 1184 122
rect 288 50 1184 122
rect 1632 50 1824 122
rect -96 122 96 986
rect 288 122 352 986
rect 1376 122 1440 986
rect 1632 122 1824 986
rect -96 986 96 1058
rect 1632 986 1824 1058
rect 288 986 352 1058
rect 416 986 1184 1058
rect 416 986 1184 1058
rect 1376 986 1440 1058
rect 1632 986 1824 1058
rect -96 1058 96 1922
rect 288 1058 352 1922
rect 1376 1058 1440 1922
rect 1632 1058 1824 1922
rect -96 1922 96 1994
rect 288 1922 1184 1994
rect 1632 1922 1824 1994
rect -96 1994 96 2080
rect 1632 1994 1824 2080
<< pcontact >>
rect 1386 338 1429 554
rect 1386 554 1429 770
rect 1386 770 1429 986
rect 1386 986 1429 1004
rect 1386 1004 1429 1022
rect 1386 1022 1429 1040
rect 1386 1040 1429 1058
rect 1386 1058 1429 1274
rect 1386 1274 1429 1490
rect 1386 1490 1429 1706
<< ptapc >>
rect -32 50 32 122
rect 1696 50 1760 122
rect -32 122 32 986
rect 1696 122 1760 986
rect -32 986 32 1058
rect 1696 986 1760 1058
rect -32 1058 32 1922
rect 1696 1058 1760 1922
rect -32 1922 32 1994
rect 1696 1922 1760 1994
<< ndcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 832 68 864 86
rect 832 86 864 104
rect 864 68 928 86
rect 864 86 928 104
rect 928 68 960 86
rect 928 86 960 104
rect 1024 68 1056 86
rect 1024 86 1056 104
rect 1056 68 1120 86
rect 1056 86 1120 104
rect 1120 68 1152 86
rect 1120 86 1152 104
rect 448 1004 480 1022
rect 448 1022 480 1040
rect 480 1004 544 1022
rect 480 1022 544 1040
rect 544 1004 576 1022
rect 544 1022 576 1040
rect 640 1004 672 1022
rect 640 1022 672 1040
rect 672 1004 736 1022
rect 672 1022 736 1040
rect 736 1004 768 1022
rect 736 1022 768 1040
rect 832 1004 864 1022
rect 832 1022 864 1040
rect 864 1004 928 1022
rect 864 1022 928 1040
rect 928 1004 960 1022
rect 928 1022 960 1040
rect 1024 1004 1056 1022
rect 1024 1022 1056 1040
rect 1056 1004 1120 1022
rect 1056 1022 1120 1040
rect 1120 1004 1152 1022
rect 1120 1022 1152 1040
rect 448 1940 480 1958
rect 448 1958 480 1976
rect 480 1940 544 1958
rect 480 1958 544 1976
rect 544 1940 576 1958
rect 544 1958 576 1976
rect 640 1940 672 1958
rect 640 1958 672 1976
rect 672 1940 736 1958
rect 672 1958 736 1976
rect 736 1940 768 1958
rect 736 1958 768 1976
rect 832 1940 864 1958
rect 832 1958 864 1976
rect 864 1940 928 1958
rect 864 1958 928 1976
rect 928 1940 960 1958
rect 928 1958 960 1976
rect 1024 1940 1056 1958
rect 1024 1958 1056 1976
rect 1056 1940 1120 1958
rect 1056 1958 1120 1976
rect 1120 1940 1152 1958
rect 1120 1958 1152 1976
<< pwell >>
rect -184 -124 1912 2168
<< labels >>
flabel locali s 1376 1058 1440 1922 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 1184 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1632 986 1824 1058 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 986 1184 1058 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1728 2030
<< end >>
