magic
tech sky130B
magscale 1 2
timestamp 1695852000
<< checkpaint >>
rect 0 0 1152 1454
<< pdiff >>
rect 416 50 608 122
rect 416 122 608 698
rect 416 698 608 770
rect 416 770 608 1346
rect 416 1346 608 1418
<< ntap >>
rect -96 -36 96 50
rect 1056 -36 1248 50
rect -96 50 96 122
rect 1056 50 1248 122
rect -96 122 96 698
rect 1056 122 1248 698
rect -96 698 96 770
rect 1056 698 1248 770
rect -96 770 96 1346
rect 1056 770 1248 1346
rect -96 1346 96 1418
rect 1056 1346 1248 1418
rect -96 1418 96 1504
rect 1056 1418 1248 1504
<< poly >>
rect 352 -18 864 32
rect 352 140 864 680
rect 352 788 864 1328
rect 352 1436 864 1486
rect 800 122 864 698
rect 800 698 864 770
rect 800 770 864 1346
<< locali >>
rect 800 770 864 1346
rect -96 -36 96 50
rect 1056 -36 1248 50
rect -96 50 96 122
rect 288 50 608 122
rect 288 50 608 122
rect 1056 50 1248 122
rect -96 122 96 698
rect 288 122 352 698
rect 800 122 864 698
rect 1056 122 1248 698
rect -96 698 96 770
rect 1056 698 1248 770
rect 288 698 352 770
rect 416 698 608 770
rect 416 698 608 770
rect 800 698 864 770
rect 1056 698 1248 770
rect -96 770 96 1346
rect 288 770 352 1346
rect 800 770 864 1346
rect 1056 770 1248 1346
rect -96 1346 96 1418
rect 288 1346 608 1418
rect 1056 1346 1248 1418
rect -96 1418 96 1504
rect 1056 1418 1248 1504
<< pcontact >>
rect 810 266 853 410
rect 810 410 853 554
rect 810 554 853 698
rect 810 698 853 716
rect 810 716 853 734
rect 810 734 853 752
rect 810 752 853 770
rect 810 770 853 914
rect 810 914 853 1058
rect 810 1058 853 1202
<< ntapc >>
rect -32 50 32 122
rect 1120 50 1184 122
rect -32 122 32 698
rect 1120 122 1184 698
rect -32 698 32 770
rect 1120 698 1184 770
rect -32 770 32 1346
rect 1120 770 1184 1346
rect -32 1346 32 1418
rect 1120 1346 1184 1418
<< pdcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 448 716 480 734
rect 448 734 480 752
rect 480 716 544 734
rect 480 734 544 752
rect 544 716 576 734
rect 544 734 576 752
rect 448 1364 480 1382
rect 448 1382 480 1400
rect 480 1364 544 1382
rect 480 1382 544 1400
rect 544 1364 576 1382
rect 544 1382 576 1400
<< nwell >>
rect -184 -124 1336 1592
<< labels >>
flabel locali s 800 770 864 1346 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 608 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1056 698 1248 770 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 698 608 770 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 1454
<< end >>
