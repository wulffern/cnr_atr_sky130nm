
*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNRATR_PCH_12C2F2_lpe.spi
#else
.include ../../../work/xsch/CNRATR_PCH_12C2F0.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-18 reltol=1e-8

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD VDD 0 dc {AVDD}
*VG 0 G dc {AVDD}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
* Passefet
XM1 OUT G VDD VDD sky130_fd_pr__pfet_01v8 L=0.252 W=11.52 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1000

* Reference
VREF VREF 0 dc 0.8
BOTA G 0 V=(1 + tanh(-1000*(v(vref) -v(out) )))/2*{AVDD}

CL OUT 0 1u

ILOAD OUT 0 pwl 0 0 1u 0 50u 0.5

BGS VGS 0 V=V(VDD)- V(G)
BIL IL 0 V=-I(VDD)



*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------


.save all
.save v(vgs)
.save i(iload)
.save v(il)


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit



optran 0 0 0 10n 10u 0

*dc VG 0.4 1.5 0.011
tran 1n 50u


write
quit
#endif

.endc

.end
