magic
tech sky130B
magscale 1 2
timestamp 1685311200
<< checkpaint >>
rect 0 0 1344 475
<< ndiff >>
rect 416 50 800 122
rect 416 122 800 208
rect 416 208 800 280
rect 416 280 800 367
rect 416 367 800 439
<< ptap >>
rect -96 -36 96 50
rect 1248 -36 1440 50
rect -96 50 96 122
rect 1248 50 1440 122
rect -96 122 96 208
rect 1248 122 1440 208
rect -96 208 96 280
rect 1248 208 1440 280
rect -96 280 96 367
rect 1248 280 1440 367
rect -96 367 96 439
rect 1248 367 1440 439
rect -96 439 96 525
rect 1248 439 1440 525
<< poly >>
rect 352 -18 1056 32
rect 352 140 1056 190
rect 352 298 1056 349
rect 352 457 1056 507
rect 992 122 1056 208
rect 992 208 1056 280
rect 992 280 1056 367
<< locali >>
rect 992 280 1056 367
rect -96 -36 96 50
rect 1248 -36 1440 50
rect -96 50 96 122
rect 288 50 800 122
rect 288 50 800 122
rect 1248 50 1440 122
rect -96 122 96 208
rect 288 122 352 208
rect 992 122 1056 208
rect 1248 122 1440 208
rect -96 208 96 280
rect 1248 208 1440 280
rect 288 208 352 280
rect 416 208 800 280
rect 416 208 800 280
rect 992 208 1056 280
rect 1248 208 1440 280
rect -96 280 96 367
rect 288 280 352 367
rect 992 280 1056 367
rect 1248 280 1440 367
rect -96 367 96 439
rect 288 367 800 439
rect 1248 367 1440 439
rect -96 439 96 525
rect 1248 439 1440 525
<< pcontact >>
rect 1002 144 1045 165
rect 1002 165 1045 187
rect 1002 187 1045 208
rect 1002 208 1045 226
rect 1002 226 1045 244
rect 1002 244 1045 262
rect 1002 262 1045 280
rect 1002 280 1045 302
rect 1002 302 1045 324
rect 1002 324 1045 345
<< ptapc >>
rect -32 50 32 122
rect 1312 50 1376 122
rect -32 122 32 208
rect 1312 122 1376 208
rect -32 208 32 280
rect 1312 208 1376 280
rect -32 280 32 367
rect 1312 280 1376 367
rect -32 367 32 439
rect 1312 367 1376 439
<< ndcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 448 226 480 244
rect 448 244 480 262
rect 480 226 544 244
rect 480 244 544 262
rect 544 226 576 244
rect 544 244 576 262
rect 640 226 672 244
rect 640 244 672 262
rect 672 226 736 244
rect 672 244 736 262
rect 736 226 768 244
rect 736 244 768 262
rect 448 385 480 403
rect 448 403 480 421
rect 480 385 544 403
rect 480 403 544 421
rect 544 385 576 403
rect 544 403 576 421
rect 640 385 672 403
rect 640 403 672 421
rect 672 385 736 403
rect 672 403 736 421
rect 736 385 768 403
rect 736 403 768 421
<< pwell >>
rect -184 -124 1528 613
<< labels >>
flabel locali s 992 280 1056 367 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 800 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1248 208 1440 280 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 208 800 280 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1344 475
<< end >>
