magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1728 1449
<< ndiff >>
rect 416 45 1184 117
rect 416 117 1184 693
rect 416 693 1184 765
rect 416 765 1184 1341
rect 416 1341 1184 1413
<< ptap >>
rect -96 -36 96 45
rect 1632 -36 1824 45
rect -96 45 96 117
rect 1632 45 1824 117
rect -96 117 96 693
rect 1632 117 1824 693
rect -96 693 96 765
rect 1632 693 1824 765
rect -96 765 96 1341
rect 1632 765 1824 1341
rect -96 1341 96 1413
rect 1632 1341 1824 1413
rect -96 1413 96 1494
rect 1632 1413 1824 1494
<< poly >>
rect 352 -18 1440 27
rect 352 135 1440 675
rect 352 783 1440 1323
rect 352 1431 1440 1476
rect 1376 117 1440 693
rect 1376 693 1440 765
rect 1376 765 1440 1341
<< locali >>
rect 1376 765 1440 1341
rect -96 -36 96 45
rect 1632 -36 1824 45
rect -96 45 96 117
rect 288 45 1184 117
rect 288 45 1184 117
rect 1632 45 1824 117
rect -96 117 96 693
rect 288 117 352 693
rect 1376 117 1440 693
rect 1632 117 1824 693
rect -96 693 96 765
rect 1632 693 1824 765
rect 288 693 352 765
rect 416 693 1184 765
rect 416 693 1184 765
rect 1376 693 1440 765
rect 1632 693 1824 765
rect -96 765 96 1341
rect 288 765 352 1341
rect 1376 765 1440 1341
rect 1632 765 1824 1341
rect -96 1341 96 1413
rect 288 1341 1184 1413
rect 1632 1341 1824 1413
rect -96 1413 96 1494
rect 1632 1413 1824 1494
<< pcontact >>
rect 1386 261 1429 405
rect 1386 405 1429 549
rect 1386 549 1429 693
rect 1386 693 1429 711
rect 1386 711 1429 729
rect 1386 729 1429 747
rect 1386 747 1429 765
rect 1386 765 1429 909
rect 1386 909 1429 1053
rect 1386 1053 1429 1197
<< ptapc >>
rect -32 45 32 117
rect 1696 45 1760 117
rect -32 117 32 693
rect 1696 117 1760 693
rect -32 693 32 765
rect 1696 693 1760 765
rect -32 765 32 1341
rect 1696 765 1760 1341
rect -32 1341 32 1413
rect 1696 1341 1760 1413
<< ndcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 832 63 864 81
rect 832 81 864 99
rect 864 63 928 81
rect 864 81 928 99
rect 928 63 960 81
rect 928 81 960 99
rect 1024 63 1056 81
rect 1024 81 1056 99
rect 1056 63 1120 81
rect 1056 81 1120 99
rect 1120 63 1152 81
rect 1120 81 1152 99
rect 448 711 480 729
rect 448 729 480 747
rect 480 711 544 729
rect 480 729 544 747
rect 544 711 576 729
rect 544 729 576 747
rect 640 711 672 729
rect 640 729 672 747
rect 672 711 736 729
rect 672 729 736 747
rect 736 711 768 729
rect 736 729 768 747
rect 832 711 864 729
rect 832 729 864 747
rect 864 711 928 729
rect 864 729 928 747
rect 928 711 960 729
rect 928 729 960 747
rect 1024 711 1056 729
rect 1024 729 1056 747
rect 1056 711 1120 729
rect 1056 729 1120 747
rect 1120 711 1152 729
rect 1120 729 1152 747
rect 448 1359 480 1377
rect 448 1377 480 1395
rect 480 1359 544 1377
rect 480 1377 544 1395
rect 544 1359 576 1377
rect 544 1377 576 1395
rect 640 1359 672 1377
rect 640 1377 672 1395
rect 672 1359 736 1377
rect 672 1377 736 1395
rect 736 1359 768 1377
rect 736 1377 768 1395
rect 832 1359 864 1377
rect 832 1377 864 1395
rect 864 1359 928 1377
rect 864 1377 928 1395
rect 928 1359 960 1377
rect 928 1377 960 1395
rect 1024 1359 1056 1377
rect 1024 1377 1056 1395
rect 1056 1359 1120 1377
rect 1056 1377 1120 1395
rect 1120 1359 1152 1377
rect 1120 1377 1152 1395
<< pwell >>
rect -184 -124 1912 1582
<< labels >>
flabel locali s 1376 765 1440 1341 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 1184 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1632 693 1824 765 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 693 1184 765 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1728 1449
<< end >>
