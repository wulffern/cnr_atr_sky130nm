magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 2112 585
<< pdiff >>
rect 416 45 1568 117
rect 416 117 1568 261
rect 416 261 1568 333
rect 416 333 1568 477
rect 416 477 1568 549
<< ntap >>
rect -96 -36 96 45
rect 2016 -36 2208 45
rect -96 45 96 117
rect 2016 45 2208 117
rect -96 117 96 261
rect 2016 117 2208 261
rect -96 261 96 333
rect 2016 261 2208 333
rect -96 333 96 477
rect 2016 333 2208 477
rect -96 477 96 549
rect 2016 477 2208 549
rect -96 549 96 630
rect 2016 549 2208 630
<< poly >>
rect 352 -18 1824 27
rect 352 135 1824 243
rect 352 351 1824 459
rect 352 567 1824 612
rect 1760 117 1824 261
rect 1760 261 1824 333
rect 1760 333 1824 477
<< locali >>
rect 1760 333 1824 477
rect -96 -36 96 45
rect 2016 -36 2208 45
rect -96 45 96 117
rect 288 45 1568 117
rect 288 45 1568 117
rect 2016 45 2208 117
rect -96 117 96 261
rect 288 117 352 261
rect 1760 117 1824 261
rect 2016 117 2208 261
rect -96 261 96 333
rect 2016 261 2208 333
rect 288 261 352 333
rect 416 261 1568 333
rect 416 261 1568 333
rect 1760 261 1824 333
rect 2016 261 2208 333
rect -96 333 96 477
rect 288 333 352 477
rect 1760 333 1824 477
rect 2016 333 2208 477
rect -96 477 96 549
rect 288 477 1568 549
rect 2016 477 2208 549
rect -96 549 96 630
rect 2016 549 2208 630
<< pcontact >>
rect 1770 153 1813 189
rect 1770 189 1813 225
rect 1770 225 1813 261
rect 1770 261 1813 279
rect 1770 279 1813 297
rect 1770 297 1813 315
rect 1770 315 1813 333
rect 1770 333 1813 369
rect 1770 369 1813 405
rect 1770 405 1813 441
<< ntapc >>
rect -32 45 32 117
rect 2080 45 2144 117
rect -32 117 32 261
rect 2080 117 2144 261
rect -32 261 32 333
rect 2080 261 2144 333
rect -32 333 32 477
rect 2080 333 2144 477
rect -32 477 32 549
rect 2080 477 2144 549
<< pdcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 832 63 864 81
rect 832 81 864 99
rect 864 63 928 81
rect 864 81 928 99
rect 928 63 960 81
rect 928 81 960 99
rect 1024 63 1056 81
rect 1024 81 1056 99
rect 1056 63 1120 81
rect 1056 81 1120 99
rect 1120 63 1152 81
rect 1120 81 1152 99
rect 1216 63 1248 81
rect 1216 81 1248 99
rect 1248 63 1312 81
rect 1248 81 1312 99
rect 1312 63 1344 81
rect 1312 81 1344 99
rect 1408 63 1440 81
rect 1408 81 1440 99
rect 1440 63 1504 81
rect 1440 81 1504 99
rect 1504 63 1536 81
rect 1504 81 1536 99
rect 448 279 480 297
rect 448 297 480 315
rect 480 279 544 297
rect 480 297 544 315
rect 544 279 576 297
rect 544 297 576 315
rect 640 279 672 297
rect 640 297 672 315
rect 672 279 736 297
rect 672 297 736 315
rect 736 279 768 297
rect 736 297 768 315
rect 832 279 864 297
rect 832 297 864 315
rect 864 279 928 297
rect 864 297 928 315
rect 928 279 960 297
rect 928 297 960 315
rect 1024 279 1056 297
rect 1024 297 1056 315
rect 1056 279 1120 297
rect 1056 297 1120 315
rect 1120 279 1152 297
rect 1120 297 1152 315
rect 1216 279 1248 297
rect 1216 297 1248 315
rect 1248 279 1312 297
rect 1248 297 1312 315
rect 1312 279 1344 297
rect 1312 297 1344 315
rect 1408 279 1440 297
rect 1408 297 1440 315
rect 1440 279 1504 297
rect 1440 297 1504 315
rect 1504 279 1536 297
rect 1504 297 1536 315
rect 448 495 480 513
rect 448 513 480 531
rect 480 495 544 513
rect 480 513 544 531
rect 544 495 576 513
rect 544 513 576 531
rect 640 495 672 513
rect 640 513 672 531
rect 672 495 736 513
rect 672 513 736 531
rect 736 495 768 513
rect 736 513 768 531
rect 832 495 864 513
rect 832 513 864 531
rect 864 495 928 513
rect 864 513 928 531
rect 928 495 960 513
rect 928 513 960 531
rect 1024 495 1056 513
rect 1024 513 1056 531
rect 1056 495 1120 513
rect 1056 513 1120 531
rect 1120 495 1152 513
rect 1120 513 1152 531
rect 1216 495 1248 513
rect 1216 513 1248 531
rect 1248 495 1312 513
rect 1248 513 1312 531
rect 1312 495 1344 513
rect 1312 513 1344 531
rect 1408 495 1440 513
rect 1408 513 1440 531
rect 1440 495 1504 513
rect 1440 513 1504 531
rect 1504 495 1536 513
rect 1504 513 1536 531
<< nwell >>
rect -184 -124 2296 718
<< labels >>
flabel locali s 1760 333 1824 477 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 1568 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 2016 261 2208 333 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 261 1568 333 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2112 585
<< end >>
