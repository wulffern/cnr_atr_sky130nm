magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1344 1449
<< pdiff >>
rect 416 45 800 117
rect 416 117 800 693
rect 416 693 800 765
rect 416 765 800 1341
rect 416 1341 800 1413
<< ntap >>
rect -96 -36 96 45
rect 1248 -36 1440 45
rect -96 45 96 117
rect 1248 45 1440 117
rect -96 117 96 693
rect 1248 117 1440 693
rect -96 693 96 765
rect 1248 693 1440 765
rect -96 765 96 1341
rect 1248 765 1440 1341
rect -96 1341 96 1413
rect 1248 1341 1440 1413
rect -96 1413 96 1494
rect 1248 1413 1440 1494
<< poly >>
rect 352 -18 1056 27
rect 352 135 1056 675
rect 352 783 1056 1323
rect 352 1431 1056 1476
rect 992 117 1056 693
rect 992 693 1056 765
rect 992 765 1056 1341
<< locali >>
rect 992 765 1056 1341
rect -96 -36 96 45
rect 1248 -36 1440 45
rect -96 45 96 117
rect 288 45 800 117
rect 288 45 800 117
rect 1248 45 1440 117
rect -96 117 96 693
rect 288 117 352 693
rect 992 117 1056 693
rect 1248 117 1440 693
rect -96 693 96 765
rect 1248 693 1440 765
rect 288 693 352 765
rect 416 693 800 765
rect 416 693 800 765
rect 992 693 1056 765
rect 1248 693 1440 765
rect -96 765 96 1341
rect 288 765 352 1341
rect 992 765 1056 1341
rect 1248 765 1440 1341
rect -96 1341 96 1413
rect 288 1341 800 1413
rect 1248 1341 1440 1413
rect -96 1413 96 1494
rect 1248 1413 1440 1494
<< pcontact >>
rect 1002 261 1045 405
rect 1002 405 1045 549
rect 1002 549 1045 693
rect 1002 693 1045 711
rect 1002 711 1045 729
rect 1002 729 1045 747
rect 1002 747 1045 765
rect 1002 765 1045 909
rect 1002 909 1045 1053
rect 1002 1053 1045 1197
<< ntapc >>
rect -32 45 32 117
rect 1312 45 1376 117
rect -32 117 32 693
rect 1312 117 1376 693
rect -32 693 32 765
rect 1312 693 1376 765
rect -32 765 32 1341
rect 1312 765 1376 1341
rect -32 1341 32 1413
rect 1312 1341 1376 1413
<< pdcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 448 711 480 729
rect 448 729 480 747
rect 480 711 544 729
rect 480 729 544 747
rect 544 711 576 729
rect 544 729 576 747
rect 640 711 672 729
rect 640 729 672 747
rect 672 711 736 729
rect 672 729 736 747
rect 736 711 768 729
rect 736 729 768 747
rect 448 1359 480 1377
rect 448 1377 480 1395
rect 480 1359 544 1377
rect 480 1377 544 1395
rect 544 1359 576 1377
rect 544 1377 576 1395
rect 640 1359 672 1377
rect 640 1377 672 1395
rect 672 1359 736 1377
rect 672 1377 736 1395
rect 736 1359 768 1377
rect 736 1377 768 1395
<< nwell >>
rect -184 -124 1528 1582
<< labels >>
flabel locali s 992 765 1056 1341 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 800 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1248 693 1440 765 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 693 800 765 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1344 1449
<< end >>
