magic
tech sky130B
magscale 1 2
timestamp 1695852000
<< checkpaint >>
rect 0 0 1152 590
<< pdiff >>
rect 416 50 608 122
rect 416 122 608 266
rect 416 266 608 338
rect 416 338 608 482
rect 416 482 608 554
<< ntap >>
rect -96 -36 96 50
rect 1056 -36 1248 50
rect -96 50 96 122
rect 1056 50 1248 122
rect -96 122 96 266
rect 1056 122 1248 266
rect -96 266 96 338
rect 1056 266 1248 338
rect -96 338 96 482
rect 1056 338 1248 482
rect -96 482 96 554
rect 1056 482 1248 554
rect -96 554 96 640
rect 1056 554 1248 640
<< poly >>
rect 352 -18 864 32
rect 352 140 864 248
rect 352 356 864 464
rect 352 572 864 622
rect 800 122 864 266
rect 800 266 864 338
rect 800 338 864 482
<< locali >>
rect 800 338 864 482
rect -96 -36 96 50
rect 1056 -36 1248 50
rect -96 50 96 122
rect 288 50 608 122
rect 288 50 608 122
rect 1056 50 1248 122
rect -96 122 96 266
rect 288 122 352 266
rect 800 122 864 266
rect 1056 122 1248 266
rect -96 266 96 338
rect 1056 266 1248 338
rect 288 266 352 338
rect 416 266 608 338
rect 416 266 608 338
rect 800 266 864 338
rect 1056 266 1248 338
rect -96 338 96 482
rect 288 338 352 482
rect 800 338 864 482
rect 1056 338 1248 482
rect -96 482 96 554
rect 288 482 608 554
rect 1056 482 1248 554
rect -96 554 96 640
rect 1056 554 1248 640
<< pcontact >>
rect 810 158 853 194
rect 810 194 853 230
rect 810 230 853 266
rect 810 266 853 284
rect 810 284 853 302
rect 810 302 853 320
rect 810 320 853 338
rect 810 338 853 374
rect 810 374 853 410
rect 810 410 853 446
<< ntapc >>
rect -32 50 32 122
rect 1120 50 1184 122
rect -32 122 32 266
rect 1120 122 1184 266
rect -32 266 32 338
rect 1120 266 1184 338
rect -32 338 32 482
rect 1120 338 1184 482
rect -32 482 32 554
rect 1120 482 1184 554
<< pdcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 448 284 480 302
rect 448 302 480 320
rect 480 284 544 302
rect 480 302 544 320
rect 544 284 576 302
rect 544 302 576 320
rect 448 500 480 518
rect 448 518 480 536
rect 480 500 544 518
rect 480 518 544 536
rect 544 500 576 518
rect 544 518 576 536
<< nwell >>
rect -184 -124 1336 728
<< labels >>
flabel locali s 800 338 864 482 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 608 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1056 266 1248 338 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 266 608 338 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 590
<< end >>
