magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1344 585
<< ndiff >>
rect 416 45 800 117
rect 416 117 800 261
rect 416 261 800 333
rect 416 333 800 477
rect 416 477 800 549
<< ptap >>
rect -96 -36 96 45
rect 1248 -36 1440 45
rect -96 45 96 117
rect 1248 45 1440 117
rect -96 117 96 261
rect 1248 117 1440 261
rect -96 261 96 333
rect 1248 261 1440 333
rect -96 333 96 477
rect 1248 333 1440 477
rect -96 477 96 549
rect 1248 477 1440 549
rect -96 549 96 630
rect 1248 549 1440 630
<< poly >>
rect 352 -18 1056 27
rect 352 135 1056 243
rect 352 351 1056 459
rect 352 567 1056 612
rect 992 117 1056 261
rect 992 261 1056 333
rect 992 333 1056 477
<< locali >>
rect 992 333 1056 477
rect -96 -36 96 45
rect 1248 -36 1440 45
rect -96 45 96 117
rect 288 45 800 117
rect 288 45 800 117
rect 1248 45 1440 117
rect -96 117 96 261
rect 288 117 352 261
rect 992 117 1056 261
rect 1248 117 1440 261
rect -96 261 96 333
rect 1248 261 1440 333
rect 288 261 352 333
rect 416 261 800 333
rect 416 261 800 333
rect 992 261 1056 333
rect 1248 261 1440 333
rect -96 333 96 477
rect 288 333 352 477
rect 992 333 1056 477
rect 1248 333 1440 477
rect -96 477 96 549
rect 288 477 800 549
rect 1248 477 1440 549
rect -96 549 96 630
rect 1248 549 1440 630
<< pcontact >>
rect 1002 153 1045 189
rect 1002 189 1045 225
rect 1002 225 1045 261
rect 1002 261 1045 279
rect 1002 279 1045 297
rect 1002 297 1045 315
rect 1002 315 1045 333
rect 1002 333 1045 369
rect 1002 369 1045 405
rect 1002 405 1045 441
<< ptapc >>
rect -32 45 32 117
rect 1312 45 1376 117
rect -32 117 32 261
rect 1312 117 1376 261
rect -32 261 32 333
rect 1312 261 1376 333
rect -32 333 32 477
rect 1312 333 1376 477
rect -32 477 32 549
rect 1312 477 1376 549
<< ndcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 448 279 480 297
rect 448 297 480 315
rect 480 279 544 297
rect 480 297 544 315
rect 544 279 576 297
rect 544 297 576 315
rect 640 279 672 297
rect 640 297 672 315
rect 672 279 736 297
rect 672 297 736 315
rect 736 279 768 297
rect 736 297 768 315
rect 448 495 480 513
rect 448 513 480 531
rect 480 495 544 513
rect 480 513 544 531
rect 544 495 576 513
rect 544 513 576 531
rect 640 495 672 513
rect 640 513 672 531
rect 672 495 736 513
rect 672 513 736 531
rect 736 495 768 513
rect 736 513 768 531
<< pwell >>
rect -184 -124 1528 718
<< labels >>
flabel locali s 992 333 1056 477 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 800 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1248 261 1440 333 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 261 800 333 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1344 585
<< end >>
