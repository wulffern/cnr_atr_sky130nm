magic
tech sky130B
magscale 1 2
timestamp 1695852000
<< checkpaint >>
rect 0 0 1344 1454
<< pdiff >>
rect 416 50 800 122
rect 416 122 800 698
rect 416 698 800 770
rect 416 770 800 1346
rect 416 1346 800 1418
<< ntap >>
rect -96 -36 96 50
rect 1248 -36 1440 50
rect -96 50 96 122
rect 1248 50 1440 122
rect -96 122 96 698
rect 1248 122 1440 698
rect -96 698 96 770
rect 1248 698 1440 770
rect -96 770 96 1346
rect 1248 770 1440 1346
rect -96 1346 96 1418
rect 1248 1346 1440 1418
rect -96 1418 96 1504
rect 1248 1418 1440 1504
<< poly >>
rect 352 -18 1056 32
rect 352 140 1056 680
rect 352 788 1056 1328
rect 352 1436 1056 1486
rect 992 122 1056 698
rect 992 698 1056 770
rect 992 770 1056 1346
<< locali >>
rect 992 770 1056 1346
rect -96 -36 96 50
rect 1248 -36 1440 50
rect -96 50 96 122
rect 288 50 800 122
rect 288 50 800 122
rect 1248 50 1440 122
rect -96 122 96 698
rect 288 122 352 698
rect 992 122 1056 698
rect 1248 122 1440 698
rect -96 698 96 770
rect 1248 698 1440 770
rect 288 698 352 770
rect 416 698 800 770
rect 416 698 800 770
rect 992 698 1056 770
rect 1248 698 1440 770
rect -96 770 96 1346
rect 288 770 352 1346
rect 992 770 1056 1346
rect 1248 770 1440 1346
rect -96 1346 96 1418
rect 288 1346 800 1418
rect 1248 1346 1440 1418
rect -96 1418 96 1504
rect 1248 1418 1440 1504
<< pcontact >>
rect 1002 266 1045 410
rect 1002 410 1045 554
rect 1002 554 1045 698
rect 1002 698 1045 716
rect 1002 716 1045 734
rect 1002 734 1045 752
rect 1002 752 1045 770
rect 1002 770 1045 914
rect 1002 914 1045 1058
rect 1002 1058 1045 1202
<< ntapc >>
rect -32 50 32 122
rect 1312 50 1376 122
rect -32 122 32 698
rect 1312 122 1376 698
rect -32 698 32 770
rect 1312 698 1376 770
rect -32 770 32 1346
rect 1312 770 1376 1346
rect -32 1346 32 1418
rect 1312 1346 1376 1418
<< pdcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 448 716 480 734
rect 448 734 480 752
rect 480 716 544 734
rect 480 734 544 752
rect 544 716 576 734
rect 544 734 576 752
rect 640 716 672 734
rect 640 734 672 752
rect 672 716 736 734
rect 672 734 736 752
rect 736 716 768 734
rect 736 734 768 752
rect 448 1364 480 1382
rect 448 1382 480 1400
rect 480 1364 544 1382
rect 480 1382 544 1400
rect 544 1364 576 1382
rect 544 1382 576 1400
rect 640 1364 672 1382
rect 640 1382 672 1400
rect 672 1364 736 1382
rect 672 1382 736 1400
rect 736 1364 768 1382
rect 736 1382 768 1400
<< nwell >>
rect -184 -124 1528 1592
<< labels >>
flabel locali s 992 770 1056 1346 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 800 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1248 698 1440 770 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 698 800 770 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1344 1454
<< end >>
