magic
tech sky130B
magscale 1 2
timestamp 1695852000
<< checkpaint >>
rect 0 0 1728 590
<< pdiff >>
rect 416 50 1184 122
rect 416 122 1184 266
rect 416 266 1184 338
rect 416 338 1184 482
rect 416 482 1184 554
<< ntap >>
rect -96 -36 96 50
rect 1632 -36 1824 50
rect -96 50 96 122
rect 1632 50 1824 122
rect -96 122 96 266
rect 1632 122 1824 266
rect -96 266 96 338
rect 1632 266 1824 338
rect -96 338 96 482
rect 1632 338 1824 482
rect -96 482 96 554
rect 1632 482 1824 554
rect -96 554 96 640
rect 1632 554 1824 640
<< poly >>
rect 352 -18 1440 32
rect 352 140 1440 248
rect 352 356 1440 464
rect 352 572 1440 622
rect 1376 122 1440 266
rect 1376 266 1440 338
rect 1376 338 1440 482
<< locali >>
rect 1376 338 1440 482
rect -96 -36 96 50
rect 1632 -36 1824 50
rect -96 50 96 122
rect 288 50 1184 122
rect 288 50 1184 122
rect 1632 50 1824 122
rect -96 122 96 266
rect 288 122 352 266
rect 1376 122 1440 266
rect 1632 122 1824 266
rect -96 266 96 338
rect 1632 266 1824 338
rect 288 266 352 338
rect 416 266 1184 338
rect 416 266 1184 338
rect 1376 266 1440 338
rect 1632 266 1824 338
rect -96 338 96 482
rect 288 338 352 482
rect 1376 338 1440 482
rect 1632 338 1824 482
rect -96 482 96 554
rect 288 482 1184 554
rect 1632 482 1824 554
rect -96 554 96 640
rect 1632 554 1824 640
<< pcontact >>
rect 1386 158 1429 194
rect 1386 194 1429 230
rect 1386 230 1429 266
rect 1386 266 1429 284
rect 1386 284 1429 302
rect 1386 302 1429 320
rect 1386 320 1429 338
rect 1386 338 1429 374
rect 1386 374 1429 410
rect 1386 410 1429 446
<< ntapc >>
rect -32 50 32 122
rect 1696 50 1760 122
rect -32 122 32 266
rect 1696 122 1760 266
rect -32 266 32 338
rect 1696 266 1760 338
rect -32 338 32 482
rect 1696 338 1760 482
rect -32 482 32 554
rect 1696 482 1760 554
<< pdcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 832 68 864 86
rect 832 86 864 104
rect 864 68 928 86
rect 864 86 928 104
rect 928 68 960 86
rect 928 86 960 104
rect 1024 68 1056 86
rect 1024 86 1056 104
rect 1056 68 1120 86
rect 1056 86 1120 104
rect 1120 68 1152 86
rect 1120 86 1152 104
rect 448 284 480 302
rect 448 302 480 320
rect 480 284 544 302
rect 480 302 544 320
rect 544 284 576 302
rect 544 302 576 320
rect 640 284 672 302
rect 640 302 672 320
rect 672 284 736 302
rect 672 302 736 320
rect 736 284 768 302
rect 736 302 768 320
rect 832 284 864 302
rect 832 302 864 320
rect 864 284 928 302
rect 864 302 928 320
rect 928 284 960 302
rect 928 302 960 320
rect 1024 284 1056 302
rect 1024 302 1056 320
rect 1056 284 1120 302
rect 1056 302 1120 320
rect 1120 284 1152 302
rect 1120 302 1152 320
rect 448 500 480 518
rect 448 518 480 536
rect 480 500 544 518
rect 480 518 544 536
rect 544 500 576 518
rect 544 518 576 536
rect 640 500 672 518
rect 640 518 672 536
rect 672 500 736 518
rect 672 518 736 536
rect 736 500 768 518
rect 736 518 768 536
rect 832 500 864 518
rect 832 518 864 536
rect 864 500 928 518
rect 864 518 928 536
rect 928 500 960 518
rect 928 518 960 536
rect 1024 500 1056 518
rect 1024 518 1056 536
rect 1056 500 1120 518
rect 1056 518 1120 536
rect 1120 500 1152 518
rect 1120 518 1152 536
<< nwell >>
rect -184 -124 1912 728
<< labels >>
flabel locali s 1376 338 1440 482 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 1184 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1632 266 1824 338 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 266 1184 338 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1728 590
<< end >>
