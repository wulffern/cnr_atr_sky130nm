magic
tech sky130B
magscale 1 2
timestamp 1685311200
<< checkpaint >>
rect 0 0 1152 878
<< ndiff >>
rect 416 50 608 122
rect 416 122 608 410
rect 416 410 608 482
rect 416 482 608 770
rect 416 770 608 842
<< ptap >>
rect -96 -36 96 50
rect 1056 -36 1248 50
rect -96 50 96 122
rect 1056 50 1248 122
rect -96 122 96 410
rect 1056 122 1248 410
rect -96 410 96 482
rect 1056 410 1248 482
rect -96 482 96 770
rect 1056 482 1248 770
rect -96 770 96 842
rect 1056 770 1248 842
rect -96 842 96 928
rect 1056 842 1248 928
<< poly >>
rect 352 -18 864 32
rect 352 140 864 392
rect 352 500 864 752
rect 352 860 864 910
rect 800 122 864 410
rect 800 410 864 482
rect 800 482 864 770
<< locali >>
rect 800 482 864 770
rect -96 -36 96 50
rect 1056 -36 1248 50
rect -96 50 96 122
rect 288 50 608 122
rect 288 50 608 122
rect 1056 50 1248 122
rect -96 122 96 410
rect 288 122 352 410
rect 800 122 864 410
rect 1056 122 1248 410
rect -96 410 96 482
rect 1056 410 1248 482
rect 288 410 352 482
rect 416 410 608 482
rect 416 410 608 482
rect 800 410 864 482
rect 1056 410 1248 482
rect -96 482 96 770
rect 288 482 352 770
rect 800 482 864 770
rect 1056 482 1248 770
rect -96 770 96 842
rect 288 770 608 842
rect 1056 770 1248 842
rect -96 842 96 928
rect 1056 842 1248 928
<< pcontact >>
rect 810 194 853 266
rect 810 266 853 338
rect 810 338 853 410
rect 810 410 853 428
rect 810 428 853 446
rect 810 446 853 464
rect 810 464 853 482
rect 810 482 853 554
rect 810 554 853 626
rect 810 626 853 698
<< ptapc >>
rect -32 50 32 122
rect 1120 50 1184 122
rect -32 122 32 410
rect 1120 122 1184 410
rect -32 410 32 482
rect 1120 410 1184 482
rect -32 482 32 770
rect 1120 482 1184 770
rect -32 770 32 842
rect 1120 770 1184 842
<< ndcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 448 428 480 446
rect 448 446 480 464
rect 480 428 544 446
rect 480 446 544 464
rect 544 428 576 446
rect 544 446 576 464
rect 448 788 480 806
rect 448 806 480 824
rect 480 788 544 806
rect 480 806 544 824
rect 544 788 576 806
rect 544 806 576 824
<< pwell >>
rect -184 -124 1336 1016
<< labels >>
flabel locali s 800 482 864 770 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 608 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1056 410 1248 482 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 410 608 482 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 878
<< end >>
