magic
tech sky130B
magscale 1 2
timestamp 1685311200
<< checkpaint >>
rect 0 0 2112 475
<< ndiff >>
rect 416 50 1568 122
rect 416 122 1568 208
rect 416 208 1568 280
rect 416 280 1568 367
rect 416 367 1568 439
<< ptap >>
rect -96 -36 96 50
rect 2016 -36 2208 50
rect -96 50 96 122
rect 2016 50 2208 122
rect -96 122 96 208
rect 2016 122 2208 208
rect -96 208 96 280
rect 2016 208 2208 280
rect -96 280 96 367
rect 2016 280 2208 367
rect -96 367 96 439
rect 2016 367 2208 439
rect -96 439 96 525
rect 2016 439 2208 525
<< poly >>
rect 352 -18 1824 32
rect 352 140 1824 190
rect 352 298 1824 349
rect 352 457 1824 507
rect 1760 122 1824 208
rect 1760 208 1824 280
rect 1760 280 1824 367
<< locali >>
rect 1760 280 1824 367
rect -96 -36 96 50
rect 2016 -36 2208 50
rect -96 50 96 122
rect 288 50 1568 122
rect 288 50 1568 122
rect 2016 50 2208 122
rect -96 122 96 208
rect 288 122 352 208
rect 1760 122 1824 208
rect 2016 122 2208 208
rect -96 208 96 280
rect 2016 208 2208 280
rect 288 208 352 280
rect 416 208 1568 280
rect 416 208 1568 280
rect 1760 208 1824 280
rect 2016 208 2208 280
rect -96 280 96 367
rect 288 280 352 367
rect 1760 280 1824 367
rect 2016 280 2208 367
rect -96 367 96 439
rect 288 367 1568 439
rect 2016 367 2208 439
rect -96 439 96 525
rect 2016 439 2208 525
<< pcontact >>
rect 1770 144 1813 165
rect 1770 165 1813 187
rect 1770 187 1813 208
rect 1770 208 1813 226
rect 1770 226 1813 244
rect 1770 244 1813 262
rect 1770 262 1813 280
rect 1770 280 1813 302
rect 1770 302 1813 324
rect 1770 324 1813 345
<< ptapc >>
rect -32 50 32 122
rect 2080 50 2144 122
rect -32 122 32 208
rect 2080 122 2144 208
rect -32 208 32 280
rect 2080 208 2144 280
rect -32 280 32 367
rect 2080 280 2144 367
rect -32 367 32 439
rect 2080 367 2144 439
<< ndcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 832 68 864 86
rect 832 86 864 104
rect 864 68 928 86
rect 864 86 928 104
rect 928 68 960 86
rect 928 86 960 104
rect 1024 68 1056 86
rect 1024 86 1056 104
rect 1056 68 1120 86
rect 1056 86 1120 104
rect 1120 68 1152 86
rect 1120 86 1152 104
rect 1216 68 1248 86
rect 1216 86 1248 104
rect 1248 68 1312 86
rect 1248 86 1312 104
rect 1312 68 1344 86
rect 1312 86 1344 104
rect 1408 68 1440 86
rect 1408 86 1440 104
rect 1440 68 1504 86
rect 1440 86 1504 104
rect 1504 68 1536 86
rect 1504 86 1536 104
rect 448 226 480 244
rect 448 244 480 262
rect 480 226 544 244
rect 480 244 544 262
rect 544 226 576 244
rect 544 244 576 262
rect 640 226 672 244
rect 640 244 672 262
rect 672 226 736 244
rect 672 244 736 262
rect 736 226 768 244
rect 736 244 768 262
rect 832 226 864 244
rect 832 244 864 262
rect 864 226 928 244
rect 864 244 928 262
rect 928 226 960 244
rect 928 244 960 262
rect 1024 226 1056 244
rect 1024 244 1056 262
rect 1056 226 1120 244
rect 1056 244 1120 262
rect 1120 226 1152 244
rect 1120 244 1152 262
rect 1216 226 1248 244
rect 1216 244 1248 262
rect 1248 226 1312 244
rect 1248 244 1312 262
rect 1312 226 1344 244
rect 1312 244 1344 262
rect 1408 226 1440 244
rect 1408 244 1440 262
rect 1440 226 1504 244
rect 1440 244 1504 262
rect 1504 226 1536 244
rect 1504 244 1536 262
rect 448 385 480 403
rect 448 403 480 421
rect 480 385 544 403
rect 480 403 544 421
rect 544 385 576 403
rect 544 403 576 421
rect 640 385 672 403
rect 640 403 672 421
rect 672 385 736 403
rect 672 403 736 421
rect 736 385 768 403
rect 736 403 768 421
rect 832 385 864 403
rect 832 403 864 421
rect 864 385 928 403
rect 864 403 928 421
rect 928 385 960 403
rect 928 403 960 421
rect 1024 385 1056 403
rect 1024 403 1056 421
rect 1056 385 1120 403
rect 1056 403 1120 421
rect 1120 385 1152 403
rect 1120 403 1152 421
rect 1216 385 1248 403
rect 1216 403 1248 421
rect 1248 385 1312 403
rect 1248 403 1312 421
rect 1312 385 1344 403
rect 1312 403 1344 421
rect 1408 385 1440 403
rect 1408 403 1440 421
rect 1440 385 1504 403
rect 1440 403 1504 421
rect 1504 385 1536 403
rect 1504 403 1536 421
<< pwell >>
rect -184 -124 2296 613
<< labels >>
flabel locali s 1760 280 1824 367 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 1568 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 2016 208 2208 280 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 208 1568 280 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2112 475
<< end >>
