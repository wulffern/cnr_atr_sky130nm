magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 2112 1449
<< ndiff >>
rect 416 45 1568 117
rect 416 117 1568 693
rect 416 693 1568 765
rect 416 765 1568 1341
rect 416 1341 1568 1413
<< ptap >>
rect -96 -36 96 45
rect 2016 -36 2208 45
rect -96 45 96 117
rect 2016 45 2208 117
rect -96 117 96 693
rect 2016 117 2208 693
rect -96 693 96 765
rect 2016 693 2208 765
rect -96 765 96 1341
rect 2016 765 2208 1341
rect -96 1341 96 1413
rect 2016 1341 2208 1413
rect -96 1413 96 1494
rect 2016 1413 2208 1494
<< poly >>
rect 352 -18 1824 27
rect 352 135 1824 675
rect 352 783 1824 1323
rect 352 1431 1824 1476
rect 1760 117 1824 693
rect 1760 693 1824 765
rect 1760 765 1824 1341
<< locali >>
rect 1760 765 1824 1341
rect -96 -36 96 45
rect 2016 -36 2208 45
rect -96 45 96 117
rect 288 45 1568 117
rect 288 45 1568 117
rect 2016 45 2208 117
rect -96 117 96 693
rect 288 117 352 693
rect 1760 117 1824 693
rect 2016 117 2208 693
rect -96 693 96 765
rect 2016 693 2208 765
rect 288 693 352 765
rect 416 693 1568 765
rect 416 693 1568 765
rect 1760 693 1824 765
rect 2016 693 2208 765
rect -96 765 96 1341
rect 288 765 352 1341
rect 1760 765 1824 1341
rect 2016 765 2208 1341
rect -96 1341 96 1413
rect 288 1341 1568 1413
rect 2016 1341 2208 1413
rect -96 1413 96 1494
rect 2016 1413 2208 1494
<< pcontact >>
rect 1770 261 1813 405
rect 1770 405 1813 549
rect 1770 549 1813 693
rect 1770 693 1813 711
rect 1770 711 1813 729
rect 1770 729 1813 747
rect 1770 747 1813 765
rect 1770 765 1813 909
rect 1770 909 1813 1053
rect 1770 1053 1813 1197
<< ptapc >>
rect -32 45 32 117
rect 2080 45 2144 117
rect -32 117 32 693
rect 2080 117 2144 693
rect -32 693 32 765
rect 2080 693 2144 765
rect -32 765 32 1341
rect 2080 765 2144 1341
rect -32 1341 32 1413
rect 2080 1341 2144 1413
<< ndcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 832 63 864 81
rect 832 81 864 99
rect 864 63 928 81
rect 864 81 928 99
rect 928 63 960 81
rect 928 81 960 99
rect 1024 63 1056 81
rect 1024 81 1056 99
rect 1056 63 1120 81
rect 1056 81 1120 99
rect 1120 63 1152 81
rect 1120 81 1152 99
rect 1216 63 1248 81
rect 1216 81 1248 99
rect 1248 63 1312 81
rect 1248 81 1312 99
rect 1312 63 1344 81
rect 1312 81 1344 99
rect 1408 63 1440 81
rect 1408 81 1440 99
rect 1440 63 1504 81
rect 1440 81 1504 99
rect 1504 63 1536 81
rect 1504 81 1536 99
rect 448 711 480 729
rect 448 729 480 747
rect 480 711 544 729
rect 480 729 544 747
rect 544 711 576 729
rect 544 729 576 747
rect 640 711 672 729
rect 640 729 672 747
rect 672 711 736 729
rect 672 729 736 747
rect 736 711 768 729
rect 736 729 768 747
rect 832 711 864 729
rect 832 729 864 747
rect 864 711 928 729
rect 864 729 928 747
rect 928 711 960 729
rect 928 729 960 747
rect 1024 711 1056 729
rect 1024 729 1056 747
rect 1056 711 1120 729
rect 1056 729 1120 747
rect 1120 711 1152 729
rect 1120 729 1152 747
rect 1216 711 1248 729
rect 1216 729 1248 747
rect 1248 711 1312 729
rect 1248 729 1312 747
rect 1312 711 1344 729
rect 1312 729 1344 747
rect 1408 711 1440 729
rect 1408 729 1440 747
rect 1440 711 1504 729
rect 1440 729 1504 747
rect 1504 711 1536 729
rect 1504 729 1536 747
rect 448 1359 480 1377
rect 448 1377 480 1395
rect 480 1359 544 1377
rect 480 1377 544 1395
rect 544 1359 576 1377
rect 544 1377 576 1395
rect 640 1359 672 1377
rect 640 1377 672 1395
rect 672 1359 736 1377
rect 672 1377 736 1395
rect 736 1359 768 1377
rect 736 1377 768 1395
rect 832 1359 864 1377
rect 832 1377 864 1395
rect 864 1359 928 1377
rect 864 1377 928 1395
rect 928 1359 960 1377
rect 928 1377 960 1395
rect 1024 1359 1056 1377
rect 1024 1377 1056 1395
rect 1056 1359 1120 1377
rect 1056 1377 1120 1395
rect 1120 1359 1152 1377
rect 1120 1377 1152 1395
rect 1216 1359 1248 1377
rect 1216 1377 1248 1395
rect 1248 1359 1312 1377
rect 1248 1377 1312 1395
rect 1312 1359 1344 1377
rect 1312 1377 1344 1395
rect 1408 1359 1440 1377
rect 1408 1377 1440 1395
rect 1440 1359 1504 1377
rect 1440 1377 1504 1395
rect 1504 1359 1536 1377
rect 1504 1377 1536 1395
<< pwell >>
rect -184 -124 2296 1582
<< labels >>
flabel locali s 1760 765 1824 1341 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 1568 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 2016 693 2208 765 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 693 1568 765 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2112 1449
<< end >>
