magic
tech sky130B
magscale 1 2
timestamp 1695852000
<< checkpaint >>
rect 0 0 1152 2030
<< pdiff >>
rect 416 50 608 122
rect 416 122 608 986
rect 416 986 608 1058
rect 416 1058 608 1922
rect 416 1922 608 1994
<< ntap >>
rect -96 -36 96 50
rect 1056 -36 1248 50
rect -96 50 96 122
rect 1056 50 1248 122
rect -96 122 96 986
rect 1056 122 1248 986
rect -96 986 96 1058
rect 1056 986 1248 1058
rect -96 1058 96 1922
rect 1056 1058 1248 1922
rect -96 1922 96 1994
rect 1056 1922 1248 1994
rect -96 1994 96 2080
rect 1056 1994 1248 2080
<< poly >>
rect 352 -18 864 32
rect 352 140 864 968
rect 352 1076 864 1904
rect 352 2012 864 2062
rect 800 122 864 986
rect 800 986 864 1058
rect 800 1058 864 1922
<< locali >>
rect 800 1058 864 1922
rect -96 -36 96 50
rect 1056 -36 1248 50
rect -96 50 96 122
rect 288 50 608 122
rect 288 50 608 122
rect 1056 50 1248 122
rect -96 122 96 986
rect 288 122 352 986
rect 800 122 864 986
rect 1056 122 1248 986
rect -96 986 96 1058
rect 1056 986 1248 1058
rect 288 986 352 1058
rect 416 986 608 1058
rect 416 986 608 1058
rect 800 986 864 1058
rect 1056 986 1248 1058
rect -96 1058 96 1922
rect 288 1058 352 1922
rect 800 1058 864 1922
rect 1056 1058 1248 1922
rect -96 1922 96 1994
rect 288 1922 608 1994
rect 1056 1922 1248 1994
rect -96 1994 96 2080
rect 1056 1994 1248 2080
<< pcontact >>
rect 810 338 853 554
rect 810 554 853 770
rect 810 770 853 986
rect 810 986 853 1004
rect 810 1004 853 1022
rect 810 1022 853 1040
rect 810 1040 853 1058
rect 810 1058 853 1274
rect 810 1274 853 1490
rect 810 1490 853 1706
<< ntapc >>
rect -32 50 32 122
rect 1120 50 1184 122
rect -32 122 32 986
rect 1120 122 1184 986
rect -32 986 32 1058
rect 1120 986 1184 1058
rect -32 1058 32 1922
rect 1120 1058 1184 1922
rect -32 1922 32 1994
rect 1120 1922 1184 1994
<< pdcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 448 1004 480 1022
rect 448 1022 480 1040
rect 480 1004 544 1022
rect 480 1022 544 1040
rect 544 1004 576 1022
rect 544 1022 576 1040
rect 448 1940 480 1958
rect 448 1958 480 1976
rect 480 1940 544 1958
rect 480 1958 544 1976
rect 544 1940 576 1958
rect 544 1958 576 1976
<< nwell >>
rect -184 -124 1336 2168
<< labels >>
flabel locali s 800 1058 864 1922 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 608 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1056 986 1248 1058 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 986 608 1058 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 2030
<< end >>
