magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1152 459
<< ndiff >>
rect 416 45 608 117
rect 416 117 608 198
rect 416 198 608 270
rect 416 270 608 351
rect 416 351 608 423
<< ptap >>
rect -96 -36 96 45
rect 1056 -36 1248 45
rect -96 45 96 117
rect 1056 45 1248 117
rect -96 117 96 198
rect 1056 117 1248 198
rect -96 198 96 270
rect 1056 198 1248 270
rect -96 270 96 351
rect 1056 270 1248 351
rect -96 351 96 423
rect 1056 351 1248 423
rect -96 423 96 504
rect 1056 423 1248 504
<< poly >>
rect 352 -18 864 27
rect 352 135 864 180
rect 352 288 864 333
rect 352 441 864 486
rect 800 117 864 198
rect 800 198 864 270
rect 800 270 864 351
<< locali >>
rect 800 270 864 351
rect -96 -36 96 45
rect 1056 -36 1248 45
rect -96 45 96 117
rect 288 45 608 117
rect 288 45 608 117
rect 1056 45 1248 117
rect -96 117 96 198
rect 288 117 352 198
rect 800 117 864 198
rect 1056 117 1248 198
rect -96 198 96 270
rect 1056 198 1248 270
rect 288 198 352 270
rect 416 198 608 270
rect 416 198 608 270
rect 800 198 864 270
rect 1056 198 1248 270
rect -96 270 96 351
rect 288 270 352 351
rect 800 270 864 351
rect 1056 270 1248 351
rect -96 351 96 423
rect 288 351 608 423
rect 1056 351 1248 423
rect -96 423 96 504
rect 1056 423 1248 504
<< pcontact >>
rect 810 137 853 157
rect 810 157 853 177
rect 810 177 853 197
rect 810 198 853 216
rect 810 216 853 234
rect 810 234 853 252
rect 810 252 853 270
rect 810 270 853 290
rect 810 290 853 310
rect 810 310 853 330
<< ptapc >>
rect -32 45 32 117
rect 1120 45 1184 117
rect -32 117 32 198
rect 1120 117 1184 198
rect -32 198 32 270
rect 1120 198 1184 270
rect -32 270 32 351
rect 1120 270 1184 351
rect -32 351 32 423
rect 1120 351 1184 423
<< ndcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 448 216 480 234
rect 448 234 480 252
rect 480 216 544 234
rect 480 234 544 252
rect 544 216 576 234
rect 544 234 576 252
rect 448 369 480 387
rect 448 387 480 405
rect 480 369 544 387
rect 480 387 544 405
rect 544 369 576 387
rect 544 387 576 405
<< pwell >>
rect -184 -124 1336 592
<< labels >>
flabel locali s 800 270 864 351 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 608 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1056 198 1248 270 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 198 608 270 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 459
<< end >>
