magic
tech sky130B
magscale 1 2
timestamp 1685311200
<< checkpaint >>
rect 0 0 1344 2030
<< ndiff >>
rect 416 50 800 122
rect 416 122 800 986
rect 416 986 800 1058
rect 416 1058 800 1922
rect 416 1922 800 1994
<< ptap >>
rect -96 -36 96 50
rect 1248 -36 1440 50
rect -96 50 96 122
rect 1248 50 1440 122
rect -96 122 96 986
rect 1248 122 1440 986
rect -96 986 96 1058
rect 1248 986 1440 1058
rect -96 1058 96 1922
rect 1248 1058 1440 1922
rect -96 1922 96 1994
rect 1248 1922 1440 1994
rect -96 1994 96 2080
rect 1248 1994 1440 2080
<< poly >>
rect 352 -18 1056 32
rect 352 140 1056 968
rect 352 1076 1056 1904
rect 352 2012 1056 2062
rect 992 122 1056 986
rect 992 986 1056 1058
rect 992 1058 1056 1922
<< locali >>
rect 992 1058 1056 1922
rect -96 -36 96 50
rect 1248 -36 1440 50
rect -96 50 96 122
rect 288 50 800 122
rect 288 50 800 122
rect 1248 50 1440 122
rect -96 122 96 986
rect 288 122 352 986
rect 992 122 1056 986
rect 1248 122 1440 986
rect -96 986 96 1058
rect 1248 986 1440 1058
rect 288 986 352 1058
rect 416 986 800 1058
rect 416 986 800 1058
rect 992 986 1056 1058
rect 1248 986 1440 1058
rect -96 1058 96 1922
rect 288 1058 352 1922
rect 992 1058 1056 1922
rect 1248 1058 1440 1922
rect -96 1922 96 1994
rect 288 1922 800 1994
rect 1248 1922 1440 1994
rect -96 1994 96 2080
rect 1248 1994 1440 2080
<< pcontact >>
rect 1002 338 1045 554
rect 1002 554 1045 770
rect 1002 770 1045 986
rect 1002 986 1045 1004
rect 1002 1004 1045 1022
rect 1002 1022 1045 1040
rect 1002 1040 1045 1058
rect 1002 1058 1045 1274
rect 1002 1274 1045 1490
rect 1002 1490 1045 1706
<< ptapc >>
rect -32 50 32 122
rect 1312 50 1376 122
rect -32 122 32 986
rect 1312 122 1376 986
rect -32 986 32 1058
rect 1312 986 1376 1058
rect -32 1058 32 1922
rect 1312 1058 1376 1922
rect -32 1922 32 1994
rect 1312 1922 1376 1994
<< ndcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 448 1004 480 1022
rect 448 1022 480 1040
rect 480 1004 544 1022
rect 480 1022 544 1040
rect 544 1004 576 1022
rect 544 1022 576 1040
rect 640 1004 672 1022
rect 640 1022 672 1040
rect 672 1004 736 1022
rect 672 1022 736 1040
rect 736 1004 768 1022
rect 736 1022 768 1040
rect 448 1940 480 1958
rect 448 1958 480 1976
rect 480 1940 544 1958
rect 480 1958 544 1976
rect 544 1940 576 1958
rect 544 1958 576 1976
rect 640 1940 672 1958
rect 640 1958 672 1976
rect 672 1940 736 1958
rect 672 1958 736 1976
rect 736 1940 768 1958
rect 736 1958 768 1976
<< pwell >>
rect -184 -124 1528 2168
<< labels >>
flabel locali s 992 1058 1056 1922 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 800 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1248 986 1440 1058 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 986 800 1058 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1344 2030
<< end >>
