magic
tech sky130B
magscale 1 2
timestamp 1685311200
<< checkpaint >>
rect 0 0 1344 878
<< pdiff >>
rect 416 50 800 122
rect 416 122 800 410
rect 416 410 800 482
rect 416 482 800 770
rect 416 770 800 842
<< ntap >>
rect -96 -36 96 50
rect 1248 -36 1440 50
rect -96 50 96 122
rect 1248 50 1440 122
rect -96 122 96 410
rect 1248 122 1440 410
rect -96 410 96 482
rect 1248 410 1440 482
rect -96 482 96 770
rect 1248 482 1440 770
rect -96 770 96 842
rect 1248 770 1440 842
rect -96 842 96 928
rect 1248 842 1440 928
<< poly >>
rect 352 -18 1056 32
rect 352 140 1056 392
rect 352 500 1056 752
rect 352 860 1056 910
rect 992 122 1056 410
rect 992 410 1056 482
rect 992 482 1056 770
<< locali >>
rect 992 482 1056 770
rect -96 -36 96 50
rect 1248 -36 1440 50
rect -96 50 96 122
rect 288 50 800 122
rect 288 50 800 122
rect 1248 50 1440 122
rect -96 122 96 410
rect 288 122 352 410
rect 992 122 1056 410
rect 1248 122 1440 410
rect -96 410 96 482
rect 1248 410 1440 482
rect 288 410 352 482
rect 416 410 800 482
rect 416 410 800 482
rect 992 410 1056 482
rect 1248 410 1440 482
rect -96 482 96 770
rect 288 482 352 770
rect 992 482 1056 770
rect 1248 482 1440 770
rect -96 770 96 842
rect 288 770 800 842
rect 1248 770 1440 842
rect -96 842 96 928
rect 1248 842 1440 928
<< pcontact >>
rect 1002 194 1045 266
rect 1002 266 1045 338
rect 1002 338 1045 410
rect 1002 410 1045 428
rect 1002 428 1045 446
rect 1002 446 1045 464
rect 1002 464 1045 482
rect 1002 482 1045 554
rect 1002 554 1045 626
rect 1002 626 1045 698
<< ntapc >>
rect -32 50 32 122
rect 1312 50 1376 122
rect -32 122 32 410
rect 1312 122 1376 410
rect -32 410 32 482
rect 1312 410 1376 482
rect -32 482 32 770
rect 1312 482 1376 770
rect -32 770 32 842
rect 1312 770 1376 842
<< pdcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 448 428 480 446
rect 448 446 480 464
rect 480 428 544 446
rect 480 446 544 464
rect 544 428 576 446
rect 544 446 576 464
rect 640 428 672 446
rect 640 446 672 464
rect 672 428 736 446
rect 672 446 736 464
rect 736 428 768 446
rect 736 446 768 464
rect 448 788 480 806
rect 448 806 480 824
rect 480 788 544 806
rect 480 806 544 824
rect 544 788 576 806
rect 544 806 576 824
rect 640 788 672 806
rect 640 806 672 824
rect 672 788 736 806
rect 672 806 736 824
rect 736 788 768 806
rect 736 806 768 824
<< nwell >>
rect -184 -124 1528 1016
<< labels >>
flabel locali s 992 482 1056 770 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 800 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1248 410 1440 482 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 410 800 482 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1344 878
<< end >>
