magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1344 2025
<< pdiff >>
rect 416 45 800 117
rect 416 117 800 981
rect 416 981 800 1053
rect 416 1053 800 1917
rect 416 1917 800 1989
<< ntap >>
rect -96 -36 96 45
rect 1248 -36 1440 45
rect -96 45 96 117
rect 1248 45 1440 117
rect -96 117 96 981
rect 1248 117 1440 981
rect -96 981 96 1053
rect 1248 981 1440 1053
rect -96 1053 96 1917
rect 1248 1053 1440 1917
rect -96 1917 96 1989
rect 1248 1917 1440 1989
rect -96 1989 96 2070
rect 1248 1989 1440 2070
<< poly >>
rect 352 -18 1056 27
rect 352 135 1056 963
rect 352 1071 1056 1899
rect 352 2007 1056 2052
rect 992 117 1056 981
rect 992 981 1056 1053
rect 992 1053 1056 1917
<< locali >>
rect 992 1053 1056 1917
rect -96 -36 96 45
rect 1248 -36 1440 45
rect -96 45 96 117
rect 288 45 800 117
rect 288 45 800 117
rect 1248 45 1440 117
rect -96 117 96 981
rect 288 117 352 981
rect 992 117 1056 981
rect 1248 117 1440 981
rect -96 981 96 1053
rect 1248 981 1440 1053
rect 288 981 352 1053
rect 416 981 800 1053
rect 416 981 800 1053
rect 992 981 1056 1053
rect 1248 981 1440 1053
rect -96 1053 96 1917
rect 288 1053 352 1917
rect 992 1053 1056 1917
rect 1248 1053 1440 1917
rect -96 1917 96 1989
rect 288 1917 800 1989
rect 1248 1917 1440 1989
rect -96 1989 96 2070
rect 1248 1989 1440 2070
<< pcontact >>
rect 1002 333 1045 549
rect 1002 549 1045 765
rect 1002 765 1045 981
rect 1002 981 1045 999
rect 1002 999 1045 1017
rect 1002 1017 1045 1035
rect 1002 1035 1045 1053
rect 1002 1053 1045 1269
rect 1002 1269 1045 1485
rect 1002 1485 1045 1701
<< ntapc >>
rect -32 45 32 117
rect 1312 45 1376 117
rect -32 117 32 981
rect 1312 117 1376 981
rect -32 981 32 1053
rect 1312 981 1376 1053
rect -32 1053 32 1917
rect 1312 1053 1376 1917
rect -32 1917 32 1989
rect 1312 1917 1376 1989
<< pdcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 448 999 480 1017
rect 448 1017 480 1035
rect 480 999 544 1017
rect 480 1017 544 1035
rect 544 999 576 1017
rect 544 1017 576 1035
rect 640 999 672 1017
rect 640 1017 672 1035
rect 672 999 736 1017
rect 672 1017 736 1035
rect 736 999 768 1017
rect 736 1017 768 1035
rect 448 1935 480 1953
rect 448 1953 480 1971
rect 480 1935 544 1953
rect 480 1953 544 1971
rect 544 1935 576 1953
rect 544 1953 576 1971
rect 640 1935 672 1953
rect 640 1953 672 1971
rect 672 1935 736 1953
rect 672 1953 736 1971
rect 736 1935 768 1953
rect 736 1953 768 1971
<< nwell >>
rect -184 -124 1528 2158
<< labels >>
flabel locali s 992 1053 1056 1917 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 800 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1248 981 1440 1053 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 981 800 1053 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1344 2025
<< end >>
