magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1344 873
<< pdiff >>
rect 416 45 800 117
rect 416 117 800 405
rect 416 405 800 477
rect 416 477 800 765
rect 416 765 800 837
<< ntap >>
rect -96 -36 96 45
rect 1248 -36 1440 45
rect -96 45 96 117
rect 1248 45 1440 117
rect -96 117 96 405
rect 1248 117 1440 405
rect -96 405 96 477
rect 1248 405 1440 477
rect -96 477 96 765
rect 1248 477 1440 765
rect -96 765 96 837
rect 1248 765 1440 837
rect -96 837 96 918
rect 1248 837 1440 918
<< poly >>
rect 352 -18 1056 27
rect 352 135 1056 387
rect 352 495 1056 747
rect 352 855 1056 900
rect 992 117 1056 405
rect 992 405 1056 477
rect 992 477 1056 765
<< locali >>
rect 992 477 1056 765
rect -96 -36 96 45
rect 1248 -36 1440 45
rect -96 45 96 117
rect 288 45 800 117
rect 288 45 800 117
rect 1248 45 1440 117
rect -96 117 96 405
rect 288 117 352 405
rect 992 117 1056 405
rect 1248 117 1440 405
rect -96 405 96 477
rect 1248 405 1440 477
rect 288 405 352 477
rect 416 405 800 477
rect 416 405 800 477
rect 992 405 1056 477
rect 1248 405 1440 477
rect -96 477 96 765
rect 288 477 352 765
rect 992 477 1056 765
rect 1248 477 1440 765
rect -96 765 96 837
rect 288 765 800 837
rect 1248 765 1440 837
rect -96 837 96 918
rect 1248 837 1440 918
<< pcontact >>
rect 1002 189 1045 261
rect 1002 261 1045 333
rect 1002 333 1045 405
rect 1002 405 1045 423
rect 1002 423 1045 441
rect 1002 441 1045 459
rect 1002 459 1045 477
rect 1002 477 1045 549
rect 1002 549 1045 621
rect 1002 621 1045 693
<< ntapc >>
rect -32 45 32 117
rect 1312 45 1376 117
rect -32 117 32 405
rect 1312 117 1376 405
rect -32 405 32 477
rect 1312 405 1376 477
rect -32 477 32 765
rect 1312 477 1376 765
rect -32 765 32 837
rect 1312 765 1376 837
<< pdcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 448 423 480 441
rect 448 441 480 459
rect 480 423 544 441
rect 480 441 544 459
rect 544 423 576 441
rect 544 441 576 459
rect 640 423 672 441
rect 640 441 672 459
rect 672 423 736 441
rect 672 441 736 459
rect 736 423 768 441
rect 736 441 768 459
rect 448 783 480 801
rect 448 801 480 819
rect 480 783 544 801
rect 480 801 544 819
rect 544 783 576 801
rect 544 801 576 819
rect 640 783 672 801
rect 640 801 672 819
rect 672 783 736 801
rect 672 801 736 819
rect 736 783 768 801
rect 736 801 768 819
<< nwell >>
rect -184 -124 1528 1006
<< labels >>
flabel locali s 992 477 1056 765 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 800 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1248 405 1440 477 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 405 800 477 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1344 873
<< end >>
