magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1728 873
<< ndiff >>
rect 416 45 1184 117
rect 416 117 1184 405
rect 416 405 1184 477
rect 416 477 1184 765
rect 416 765 1184 837
<< ptap >>
rect -96 -36 96 45
rect 1632 -36 1824 45
rect -96 45 96 117
rect 1632 45 1824 117
rect -96 117 96 405
rect 1632 117 1824 405
rect -96 405 96 477
rect 1632 405 1824 477
rect -96 477 96 765
rect 1632 477 1824 765
rect -96 765 96 837
rect 1632 765 1824 837
rect -96 837 96 918
rect 1632 837 1824 918
<< poly >>
rect 352 -18 1440 27
rect 352 135 1440 387
rect 352 495 1440 747
rect 352 855 1440 900
rect 1376 117 1440 405
rect 1376 405 1440 477
rect 1376 477 1440 765
<< locali >>
rect 1376 477 1440 765
rect -96 -36 96 45
rect 1632 -36 1824 45
rect -96 45 96 117
rect 288 45 1184 117
rect 288 45 1184 117
rect 1632 45 1824 117
rect -96 117 96 405
rect 288 117 352 405
rect 1376 117 1440 405
rect 1632 117 1824 405
rect -96 405 96 477
rect 1632 405 1824 477
rect 288 405 352 477
rect 416 405 1184 477
rect 416 405 1184 477
rect 1376 405 1440 477
rect 1632 405 1824 477
rect -96 477 96 765
rect 288 477 352 765
rect 1376 477 1440 765
rect 1632 477 1824 765
rect -96 765 96 837
rect 288 765 1184 837
rect 1632 765 1824 837
rect -96 837 96 918
rect 1632 837 1824 918
<< pcontact >>
rect 1386 189 1429 261
rect 1386 261 1429 333
rect 1386 333 1429 405
rect 1386 405 1429 423
rect 1386 423 1429 441
rect 1386 441 1429 459
rect 1386 459 1429 477
rect 1386 477 1429 549
rect 1386 549 1429 621
rect 1386 621 1429 693
<< ptapc >>
rect -32 45 32 117
rect 1696 45 1760 117
rect -32 117 32 405
rect 1696 117 1760 405
rect -32 405 32 477
rect 1696 405 1760 477
rect -32 477 32 765
rect 1696 477 1760 765
rect -32 765 32 837
rect 1696 765 1760 837
<< ndcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 832 63 864 81
rect 832 81 864 99
rect 864 63 928 81
rect 864 81 928 99
rect 928 63 960 81
rect 928 81 960 99
rect 1024 63 1056 81
rect 1024 81 1056 99
rect 1056 63 1120 81
rect 1056 81 1120 99
rect 1120 63 1152 81
rect 1120 81 1152 99
rect 448 423 480 441
rect 448 441 480 459
rect 480 423 544 441
rect 480 441 544 459
rect 544 423 576 441
rect 544 441 576 459
rect 640 423 672 441
rect 640 441 672 459
rect 672 423 736 441
rect 672 441 736 459
rect 736 423 768 441
rect 736 441 768 459
rect 832 423 864 441
rect 832 441 864 459
rect 864 423 928 441
rect 864 441 928 459
rect 928 423 960 441
rect 928 441 960 459
rect 1024 423 1056 441
rect 1024 441 1056 459
rect 1056 423 1120 441
rect 1056 441 1120 459
rect 1120 423 1152 441
rect 1120 441 1152 459
rect 448 783 480 801
rect 448 801 480 819
rect 480 783 544 801
rect 480 801 544 819
rect 544 783 576 801
rect 544 801 576 819
rect 640 783 672 801
rect 640 801 672 819
rect 672 783 736 801
rect 672 801 736 819
rect 736 783 768 801
rect 736 801 768 819
rect 832 783 864 801
rect 832 801 864 819
rect 864 783 928 801
rect 864 801 928 819
rect 928 783 960 801
rect 928 801 960 819
rect 1024 783 1056 801
rect 1024 801 1056 819
rect 1056 783 1120 801
rect 1056 801 1120 819
rect 1120 783 1152 801
rect 1120 801 1152 819
<< pwell >>
rect -184 -124 1912 1006
<< labels >>
flabel locali s 1376 477 1440 765 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 1184 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1632 405 1824 477 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 405 1184 477 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1728 873
<< end >>
