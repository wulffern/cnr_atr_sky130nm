magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1152 1449
<< pdiff >>
rect 416 45 608 117
rect 416 117 608 693
rect 416 693 608 765
rect 416 765 608 1341
rect 416 1341 608 1413
<< ntap >>
rect -96 -36 96 45
rect 1056 -36 1248 45
rect -96 45 96 117
rect 1056 45 1248 117
rect -96 117 96 693
rect 1056 117 1248 693
rect -96 693 96 765
rect 1056 693 1248 765
rect -96 765 96 1341
rect 1056 765 1248 1341
rect -96 1341 96 1413
rect 1056 1341 1248 1413
rect -96 1413 96 1494
rect 1056 1413 1248 1494
<< poly >>
rect 352 -18 864 27
rect 352 135 864 675
rect 352 783 864 1323
rect 352 1431 864 1476
rect 800 117 864 693
rect 800 693 864 765
rect 800 765 864 1341
<< locali >>
rect 800 765 864 1341
rect -96 -36 96 45
rect 1056 -36 1248 45
rect -96 45 96 117
rect 288 45 608 117
rect 288 45 608 117
rect 1056 45 1248 117
rect -96 117 96 693
rect 288 117 352 693
rect 800 117 864 693
rect 1056 117 1248 693
rect -96 693 96 765
rect 1056 693 1248 765
rect 288 693 352 765
rect 416 693 608 765
rect 416 693 608 765
rect 800 693 864 765
rect 1056 693 1248 765
rect -96 765 96 1341
rect 288 765 352 1341
rect 800 765 864 1341
rect 1056 765 1248 1341
rect -96 1341 96 1413
rect 288 1341 608 1413
rect 1056 1341 1248 1413
rect -96 1413 96 1494
rect 1056 1413 1248 1494
<< pcontact >>
rect 810 261 853 405
rect 810 405 853 549
rect 810 549 853 693
rect 810 693 853 711
rect 810 711 853 729
rect 810 729 853 747
rect 810 747 853 765
rect 810 765 853 909
rect 810 909 853 1053
rect 810 1053 853 1197
<< ntapc >>
rect -32 45 32 117
rect 1120 45 1184 117
rect -32 117 32 693
rect 1120 117 1184 693
rect -32 693 32 765
rect 1120 693 1184 765
rect -32 765 32 1341
rect 1120 765 1184 1341
rect -32 1341 32 1413
rect 1120 1341 1184 1413
<< pdcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 448 711 480 729
rect 448 729 480 747
rect 480 711 544 729
rect 480 729 544 747
rect 544 711 576 729
rect 544 729 576 747
rect 448 1359 480 1377
rect 448 1377 480 1395
rect 480 1359 544 1377
rect 480 1377 544 1395
rect 544 1359 576 1377
rect 544 1377 576 1395
<< nwell >>
rect -184 -124 1336 1582
<< labels >>
flabel locali s 800 765 864 1341 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 608 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1056 693 1248 765 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 693 608 765 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 1449
<< end >>
