magic
tech sky130B
magscale 1 2
timestamp 1685311200
<< checkpaint >>
rect 0 0 2112 2030
<< ndiff >>
rect 416 50 1568 122
rect 416 122 1568 986
rect 416 986 1568 1058
rect 416 1058 1568 1922
rect 416 1922 1568 1994
<< ptap >>
rect -96 -36 96 50
rect 2016 -36 2208 50
rect -96 50 96 122
rect 2016 50 2208 122
rect -96 122 96 986
rect 2016 122 2208 986
rect -96 986 96 1058
rect 2016 986 2208 1058
rect -96 1058 96 1922
rect 2016 1058 2208 1922
rect -96 1922 96 1994
rect 2016 1922 2208 1994
rect -96 1994 96 2080
rect 2016 1994 2208 2080
<< poly >>
rect 352 -18 1824 32
rect 352 140 1824 968
rect 352 1076 1824 1904
rect 352 2012 1824 2062
rect 1760 122 1824 986
rect 1760 986 1824 1058
rect 1760 1058 1824 1922
<< locali >>
rect 1760 1058 1824 1922
rect -96 -36 96 50
rect 2016 -36 2208 50
rect -96 50 96 122
rect 288 50 1568 122
rect 288 50 1568 122
rect 2016 50 2208 122
rect -96 122 96 986
rect 288 122 352 986
rect 1760 122 1824 986
rect 2016 122 2208 986
rect -96 986 96 1058
rect 2016 986 2208 1058
rect 288 986 352 1058
rect 416 986 1568 1058
rect 416 986 1568 1058
rect 1760 986 1824 1058
rect 2016 986 2208 1058
rect -96 1058 96 1922
rect 288 1058 352 1922
rect 1760 1058 1824 1922
rect 2016 1058 2208 1922
rect -96 1922 96 1994
rect 288 1922 1568 1994
rect 2016 1922 2208 1994
rect -96 1994 96 2080
rect 2016 1994 2208 2080
<< pcontact >>
rect 1770 338 1813 554
rect 1770 554 1813 770
rect 1770 770 1813 986
rect 1770 986 1813 1004
rect 1770 1004 1813 1022
rect 1770 1022 1813 1040
rect 1770 1040 1813 1058
rect 1770 1058 1813 1274
rect 1770 1274 1813 1490
rect 1770 1490 1813 1706
<< ptapc >>
rect -32 50 32 122
rect 2080 50 2144 122
rect -32 122 32 986
rect 2080 122 2144 986
rect -32 986 32 1058
rect 2080 986 2144 1058
rect -32 1058 32 1922
rect 2080 1058 2144 1922
rect -32 1922 32 1994
rect 2080 1922 2144 1994
<< ndcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 832 68 864 86
rect 832 86 864 104
rect 864 68 928 86
rect 864 86 928 104
rect 928 68 960 86
rect 928 86 960 104
rect 1024 68 1056 86
rect 1024 86 1056 104
rect 1056 68 1120 86
rect 1056 86 1120 104
rect 1120 68 1152 86
rect 1120 86 1152 104
rect 1216 68 1248 86
rect 1216 86 1248 104
rect 1248 68 1312 86
rect 1248 86 1312 104
rect 1312 68 1344 86
rect 1312 86 1344 104
rect 1408 68 1440 86
rect 1408 86 1440 104
rect 1440 68 1504 86
rect 1440 86 1504 104
rect 1504 68 1536 86
rect 1504 86 1536 104
rect 448 1004 480 1022
rect 448 1022 480 1040
rect 480 1004 544 1022
rect 480 1022 544 1040
rect 544 1004 576 1022
rect 544 1022 576 1040
rect 640 1004 672 1022
rect 640 1022 672 1040
rect 672 1004 736 1022
rect 672 1022 736 1040
rect 736 1004 768 1022
rect 736 1022 768 1040
rect 832 1004 864 1022
rect 832 1022 864 1040
rect 864 1004 928 1022
rect 864 1022 928 1040
rect 928 1004 960 1022
rect 928 1022 960 1040
rect 1024 1004 1056 1022
rect 1024 1022 1056 1040
rect 1056 1004 1120 1022
rect 1056 1022 1120 1040
rect 1120 1004 1152 1022
rect 1120 1022 1152 1040
rect 1216 1004 1248 1022
rect 1216 1022 1248 1040
rect 1248 1004 1312 1022
rect 1248 1022 1312 1040
rect 1312 1004 1344 1022
rect 1312 1022 1344 1040
rect 1408 1004 1440 1022
rect 1408 1022 1440 1040
rect 1440 1004 1504 1022
rect 1440 1022 1504 1040
rect 1504 1004 1536 1022
rect 1504 1022 1536 1040
rect 448 1940 480 1958
rect 448 1958 480 1976
rect 480 1940 544 1958
rect 480 1958 544 1976
rect 544 1940 576 1958
rect 544 1958 576 1976
rect 640 1940 672 1958
rect 640 1958 672 1976
rect 672 1940 736 1958
rect 672 1958 736 1976
rect 736 1940 768 1958
rect 736 1958 768 1976
rect 832 1940 864 1958
rect 832 1958 864 1976
rect 864 1940 928 1958
rect 864 1958 928 1976
rect 928 1940 960 1958
rect 928 1958 960 1976
rect 1024 1940 1056 1958
rect 1024 1958 1056 1976
rect 1056 1940 1120 1958
rect 1056 1958 1120 1976
rect 1120 1940 1152 1958
rect 1120 1958 1152 1976
rect 1216 1940 1248 1958
rect 1216 1958 1248 1976
rect 1248 1940 1312 1958
rect 1248 1958 1312 1976
rect 1312 1940 1344 1958
rect 1312 1958 1344 1976
rect 1408 1940 1440 1958
rect 1408 1958 1440 1976
rect 1440 1940 1504 1958
rect 1440 1958 1504 1976
rect 1504 1940 1536 1958
rect 1504 1958 1536 1976
<< pwell >>
rect -184 -124 2296 2168
<< labels >>
flabel locali s 1760 1058 1824 1922 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 1568 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 2016 986 2208 1058 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 986 1568 1058 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2112 2030
<< end >>
