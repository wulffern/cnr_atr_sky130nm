magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1152 873
<< ndiff >>
rect 416 45 608 117
rect 416 117 608 405
rect 416 405 608 477
rect 416 477 608 765
rect 416 765 608 837
<< ptap >>
rect -96 -36 96 45
rect 1056 -36 1248 45
rect -96 45 96 117
rect 1056 45 1248 117
rect -96 117 96 405
rect 1056 117 1248 405
rect -96 405 96 477
rect 1056 405 1248 477
rect -96 477 96 765
rect 1056 477 1248 765
rect -96 765 96 837
rect 1056 765 1248 837
rect -96 837 96 918
rect 1056 837 1248 918
<< poly >>
rect 352 -18 864 27
rect 352 135 864 387
rect 352 495 864 747
rect 352 855 864 900
rect 800 117 864 405
rect 800 405 864 477
rect 800 477 864 765
<< locali >>
rect 800 477 864 765
rect -96 -36 96 45
rect 1056 -36 1248 45
rect -96 45 96 117
rect 288 45 608 117
rect 288 45 608 117
rect 1056 45 1248 117
rect -96 117 96 405
rect 288 117 352 405
rect 800 117 864 405
rect 1056 117 1248 405
rect -96 405 96 477
rect 1056 405 1248 477
rect 288 405 352 477
rect 416 405 608 477
rect 416 405 608 477
rect 800 405 864 477
rect 1056 405 1248 477
rect -96 477 96 765
rect 288 477 352 765
rect 800 477 864 765
rect 1056 477 1248 765
rect -96 765 96 837
rect 288 765 608 837
rect 1056 765 1248 837
rect -96 837 96 918
rect 1056 837 1248 918
<< pcontact >>
rect 810 189 853 261
rect 810 261 853 333
rect 810 333 853 405
rect 810 405 853 423
rect 810 423 853 441
rect 810 441 853 459
rect 810 459 853 477
rect 810 477 853 549
rect 810 549 853 621
rect 810 621 853 693
<< ptapc >>
rect -32 45 32 117
rect 1120 45 1184 117
rect -32 117 32 405
rect 1120 117 1184 405
rect -32 405 32 477
rect 1120 405 1184 477
rect -32 477 32 765
rect 1120 477 1184 765
rect -32 765 32 837
rect 1120 765 1184 837
<< ndcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 448 423 480 441
rect 448 441 480 459
rect 480 423 544 441
rect 480 441 544 459
rect 544 423 576 441
rect 544 441 576 459
rect 448 783 480 801
rect 448 801 480 819
rect 480 783 544 801
rect 480 801 544 819
rect 544 783 576 801
rect 544 801 576 819
<< pwell >>
rect -184 -124 1336 1006
<< labels >>
flabel locali s 800 477 864 765 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 608 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1056 405 1248 477 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 405 608 477 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 873
<< end >>
