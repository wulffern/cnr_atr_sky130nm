magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1728 585
<< ndiff >>
rect 416 45 1184 117
rect 416 117 1184 261
rect 416 261 1184 333
rect 416 333 1184 477
rect 416 477 1184 549
<< ptap >>
rect -96 -36 96 45
rect 1632 -36 1824 45
rect -96 45 96 117
rect 1632 45 1824 117
rect -96 117 96 261
rect 1632 117 1824 261
rect -96 261 96 333
rect 1632 261 1824 333
rect -96 333 96 477
rect 1632 333 1824 477
rect -96 477 96 549
rect 1632 477 1824 549
rect -96 549 96 630
rect 1632 549 1824 630
<< poly >>
rect 352 -18 1440 27
rect 352 135 1440 243
rect 352 351 1440 459
rect 352 567 1440 612
rect 1376 117 1440 261
rect 1376 261 1440 333
rect 1376 333 1440 477
<< locali >>
rect 1376 333 1440 477
rect -96 -36 96 45
rect 1632 -36 1824 45
rect -96 45 96 117
rect 288 45 1184 117
rect 288 45 1184 117
rect 1632 45 1824 117
rect -96 117 96 261
rect 288 117 352 261
rect 1376 117 1440 261
rect 1632 117 1824 261
rect -96 261 96 333
rect 1632 261 1824 333
rect 288 261 352 333
rect 416 261 1184 333
rect 416 261 1184 333
rect 1376 261 1440 333
rect 1632 261 1824 333
rect -96 333 96 477
rect 288 333 352 477
rect 1376 333 1440 477
rect 1632 333 1824 477
rect -96 477 96 549
rect 288 477 1184 549
rect 1632 477 1824 549
rect -96 549 96 630
rect 1632 549 1824 630
<< pcontact >>
rect 1386 153 1429 189
rect 1386 189 1429 225
rect 1386 225 1429 261
rect 1386 261 1429 279
rect 1386 279 1429 297
rect 1386 297 1429 315
rect 1386 315 1429 333
rect 1386 333 1429 369
rect 1386 369 1429 405
rect 1386 405 1429 441
<< ptapc >>
rect -32 45 32 117
rect 1696 45 1760 117
rect -32 117 32 261
rect 1696 117 1760 261
rect -32 261 32 333
rect 1696 261 1760 333
rect -32 333 32 477
rect 1696 333 1760 477
rect -32 477 32 549
rect 1696 477 1760 549
<< ndcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 832 63 864 81
rect 832 81 864 99
rect 864 63 928 81
rect 864 81 928 99
rect 928 63 960 81
rect 928 81 960 99
rect 1024 63 1056 81
rect 1024 81 1056 99
rect 1056 63 1120 81
rect 1056 81 1120 99
rect 1120 63 1152 81
rect 1120 81 1152 99
rect 448 279 480 297
rect 448 297 480 315
rect 480 279 544 297
rect 480 297 544 315
rect 544 279 576 297
rect 544 297 576 315
rect 640 279 672 297
rect 640 297 672 315
rect 672 279 736 297
rect 672 297 736 315
rect 736 279 768 297
rect 736 297 768 315
rect 832 279 864 297
rect 832 297 864 315
rect 864 279 928 297
rect 864 297 928 315
rect 928 279 960 297
rect 928 297 960 315
rect 1024 279 1056 297
rect 1024 297 1056 315
rect 1056 279 1120 297
rect 1056 297 1120 315
rect 1120 279 1152 297
rect 1120 297 1152 315
rect 448 495 480 513
rect 448 513 480 531
rect 480 495 544 513
rect 480 513 544 531
rect 544 495 576 513
rect 544 513 576 531
rect 640 495 672 513
rect 640 513 672 531
rect 672 495 736 513
rect 672 513 736 531
rect 736 495 768 513
rect 736 513 768 531
rect 832 495 864 513
rect 832 513 864 531
rect 864 495 928 513
rect 864 513 928 531
rect 928 495 960 513
rect 928 513 960 531
rect 1024 495 1056 513
rect 1024 513 1056 531
rect 1056 495 1120 513
rect 1056 513 1120 531
rect 1120 495 1152 513
rect 1120 513 1152 531
<< pwell >>
rect -184 -124 1912 718
<< labels >>
flabel locali s 1376 333 1440 477 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 1184 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1632 261 1824 333 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 261 1184 333 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1728 585
<< end >>
