magic
tech sky130B
magscale 1 2
timestamp 1695852000
<< checkpaint >>
rect 0 0 2112 878
<< pdiff >>
rect 416 50 1568 122
rect 416 122 1568 410
rect 416 410 1568 482
rect 416 482 1568 770
rect 416 770 1568 842
<< ntap >>
rect -96 -36 96 50
rect 2016 -36 2208 50
rect -96 50 96 122
rect 2016 50 2208 122
rect -96 122 96 410
rect 2016 122 2208 410
rect -96 410 96 482
rect 2016 410 2208 482
rect -96 482 96 770
rect 2016 482 2208 770
rect -96 770 96 842
rect 2016 770 2208 842
rect -96 842 96 928
rect 2016 842 2208 928
<< poly >>
rect 352 -18 1824 32
rect 352 140 1824 392
rect 352 500 1824 752
rect 352 860 1824 910
rect 1760 122 1824 410
rect 1760 410 1824 482
rect 1760 482 1824 770
<< locali >>
rect 1760 482 1824 770
rect -96 -36 96 50
rect 2016 -36 2208 50
rect -96 50 96 122
rect 288 50 1568 122
rect 288 50 1568 122
rect 2016 50 2208 122
rect -96 122 96 410
rect 288 122 352 410
rect 1760 122 1824 410
rect 2016 122 2208 410
rect -96 410 96 482
rect 2016 410 2208 482
rect 288 410 352 482
rect 416 410 1568 482
rect 416 410 1568 482
rect 1760 410 1824 482
rect 2016 410 2208 482
rect -96 482 96 770
rect 288 482 352 770
rect 1760 482 1824 770
rect 2016 482 2208 770
rect -96 770 96 842
rect 288 770 1568 842
rect 2016 770 2208 842
rect -96 842 96 928
rect 2016 842 2208 928
<< pcontact >>
rect 1770 194 1813 266
rect 1770 266 1813 338
rect 1770 338 1813 410
rect 1770 410 1813 428
rect 1770 428 1813 446
rect 1770 446 1813 464
rect 1770 464 1813 482
rect 1770 482 1813 554
rect 1770 554 1813 626
rect 1770 626 1813 698
<< ntapc >>
rect -32 50 32 122
rect 2080 50 2144 122
rect -32 122 32 410
rect 2080 122 2144 410
rect -32 410 32 482
rect 2080 410 2144 482
rect -32 482 32 770
rect 2080 482 2144 770
rect -32 770 32 842
rect 2080 770 2144 842
<< pdcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 832 68 864 86
rect 832 86 864 104
rect 864 68 928 86
rect 864 86 928 104
rect 928 68 960 86
rect 928 86 960 104
rect 1024 68 1056 86
rect 1024 86 1056 104
rect 1056 68 1120 86
rect 1056 86 1120 104
rect 1120 68 1152 86
rect 1120 86 1152 104
rect 1216 68 1248 86
rect 1216 86 1248 104
rect 1248 68 1312 86
rect 1248 86 1312 104
rect 1312 68 1344 86
rect 1312 86 1344 104
rect 1408 68 1440 86
rect 1408 86 1440 104
rect 1440 68 1504 86
rect 1440 86 1504 104
rect 1504 68 1536 86
rect 1504 86 1536 104
rect 448 428 480 446
rect 448 446 480 464
rect 480 428 544 446
rect 480 446 544 464
rect 544 428 576 446
rect 544 446 576 464
rect 640 428 672 446
rect 640 446 672 464
rect 672 428 736 446
rect 672 446 736 464
rect 736 428 768 446
rect 736 446 768 464
rect 832 428 864 446
rect 832 446 864 464
rect 864 428 928 446
rect 864 446 928 464
rect 928 428 960 446
rect 928 446 960 464
rect 1024 428 1056 446
rect 1024 446 1056 464
rect 1056 428 1120 446
rect 1056 446 1120 464
rect 1120 428 1152 446
rect 1120 446 1152 464
rect 1216 428 1248 446
rect 1216 446 1248 464
rect 1248 428 1312 446
rect 1248 446 1312 464
rect 1312 428 1344 446
rect 1312 446 1344 464
rect 1408 428 1440 446
rect 1408 446 1440 464
rect 1440 428 1504 446
rect 1440 446 1504 464
rect 1504 428 1536 446
rect 1504 446 1536 464
rect 448 788 480 806
rect 448 806 480 824
rect 480 788 544 806
rect 480 806 544 824
rect 544 788 576 806
rect 544 806 576 824
rect 640 788 672 806
rect 640 806 672 824
rect 672 788 736 806
rect 672 806 736 824
rect 736 788 768 806
rect 736 806 768 824
rect 832 788 864 806
rect 832 806 864 824
rect 864 788 928 806
rect 864 806 928 824
rect 928 788 960 806
rect 928 806 960 824
rect 1024 788 1056 806
rect 1024 806 1056 824
rect 1056 788 1120 806
rect 1056 806 1120 824
rect 1120 788 1152 806
rect 1120 806 1152 824
rect 1216 788 1248 806
rect 1216 806 1248 824
rect 1248 788 1312 806
rect 1248 806 1312 824
rect 1312 788 1344 806
rect 1312 806 1344 824
rect 1408 788 1440 806
rect 1408 806 1440 824
rect 1440 788 1504 806
rect 1440 806 1504 824
rect 1504 788 1536 806
rect 1504 806 1536 824
<< nwell >>
rect -184 -124 2296 1016
<< labels >>
flabel locali s 1760 482 1824 770 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 1568 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 2016 410 2208 482 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 410 1568 482 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2112 878
<< end >>
