magic
tech sky130B
magscale 1 2
timestamp 1695852000
<< checkpaint >>
rect 0 0 1344 590
<< pdiff >>
rect 416 50 800 122
rect 416 122 800 266
rect 416 266 800 338
rect 416 338 800 482
rect 416 482 800 554
<< ntap >>
rect -96 -36 96 50
rect 1248 -36 1440 50
rect -96 50 96 122
rect 1248 50 1440 122
rect -96 122 96 266
rect 1248 122 1440 266
rect -96 266 96 338
rect 1248 266 1440 338
rect -96 338 96 482
rect 1248 338 1440 482
rect -96 482 96 554
rect 1248 482 1440 554
rect -96 554 96 640
rect 1248 554 1440 640
<< poly >>
rect 352 -18 1056 32
rect 352 140 1056 248
rect 352 356 1056 464
rect 352 572 1056 622
rect 992 122 1056 266
rect 992 266 1056 338
rect 992 338 1056 482
<< locali >>
rect 992 338 1056 482
rect -96 -36 96 50
rect 1248 -36 1440 50
rect -96 50 96 122
rect 288 50 800 122
rect 288 50 800 122
rect 1248 50 1440 122
rect -96 122 96 266
rect 288 122 352 266
rect 992 122 1056 266
rect 1248 122 1440 266
rect -96 266 96 338
rect 1248 266 1440 338
rect 288 266 352 338
rect 416 266 800 338
rect 416 266 800 338
rect 992 266 1056 338
rect 1248 266 1440 338
rect -96 338 96 482
rect 288 338 352 482
rect 992 338 1056 482
rect 1248 338 1440 482
rect -96 482 96 554
rect 288 482 800 554
rect 1248 482 1440 554
rect -96 554 96 640
rect 1248 554 1440 640
<< pcontact >>
rect 1002 158 1045 194
rect 1002 194 1045 230
rect 1002 230 1045 266
rect 1002 266 1045 284
rect 1002 284 1045 302
rect 1002 302 1045 320
rect 1002 320 1045 338
rect 1002 338 1045 374
rect 1002 374 1045 410
rect 1002 410 1045 446
<< ntapc >>
rect -32 50 32 122
rect 1312 50 1376 122
rect -32 122 32 266
rect 1312 122 1376 266
rect -32 266 32 338
rect 1312 266 1376 338
rect -32 338 32 482
rect 1312 338 1376 482
rect -32 482 32 554
rect 1312 482 1376 554
<< pdcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 448 284 480 302
rect 448 302 480 320
rect 480 284 544 302
rect 480 302 544 320
rect 544 284 576 302
rect 544 302 576 320
rect 640 284 672 302
rect 640 302 672 320
rect 672 284 736 302
rect 672 302 736 320
rect 736 284 768 302
rect 736 302 768 320
rect 448 500 480 518
rect 448 518 480 536
rect 480 500 544 518
rect 480 518 544 536
rect 544 500 576 518
rect 544 518 576 536
rect 640 500 672 518
rect 640 518 672 536
rect 672 500 736 518
rect 672 518 736 536
rect 736 500 768 518
rect 736 518 768 536
<< nwell >>
rect -184 -124 1528 728
<< labels >>
flabel locali s 992 338 1056 482 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 800 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1248 266 1440 338 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 266 800 338 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1344 590
<< end >>
