magic
tech sky130B
magscale 1 2
timestamp 1695852000
<< checkpaint >>
rect 0 0 2112 590
<< pdiff >>
rect 416 50 1568 122
rect 416 122 1568 266
rect 416 266 1568 338
rect 416 338 1568 482
rect 416 482 1568 554
<< ntap >>
rect -96 -36 96 50
rect 2016 -36 2208 50
rect -96 50 96 122
rect 2016 50 2208 122
rect -96 122 96 266
rect 2016 122 2208 266
rect -96 266 96 338
rect 2016 266 2208 338
rect -96 338 96 482
rect 2016 338 2208 482
rect -96 482 96 554
rect 2016 482 2208 554
rect -96 554 96 640
rect 2016 554 2208 640
<< poly >>
rect 352 -18 1824 32
rect 352 140 1824 248
rect 352 356 1824 464
rect 352 572 1824 622
rect 1760 122 1824 266
rect 1760 266 1824 338
rect 1760 338 1824 482
<< locali >>
rect 1760 338 1824 482
rect -96 -36 96 50
rect 2016 -36 2208 50
rect -96 50 96 122
rect 288 50 1568 122
rect 288 50 1568 122
rect 2016 50 2208 122
rect -96 122 96 266
rect 288 122 352 266
rect 1760 122 1824 266
rect 2016 122 2208 266
rect -96 266 96 338
rect 2016 266 2208 338
rect 288 266 352 338
rect 416 266 1568 338
rect 416 266 1568 338
rect 1760 266 1824 338
rect 2016 266 2208 338
rect -96 338 96 482
rect 288 338 352 482
rect 1760 338 1824 482
rect 2016 338 2208 482
rect -96 482 96 554
rect 288 482 1568 554
rect 2016 482 2208 554
rect -96 554 96 640
rect 2016 554 2208 640
<< pcontact >>
rect 1770 158 1813 194
rect 1770 194 1813 230
rect 1770 230 1813 266
rect 1770 266 1813 284
rect 1770 284 1813 302
rect 1770 302 1813 320
rect 1770 320 1813 338
rect 1770 338 1813 374
rect 1770 374 1813 410
rect 1770 410 1813 446
<< ntapc >>
rect -32 50 32 122
rect 2080 50 2144 122
rect -32 122 32 266
rect 2080 122 2144 266
rect -32 266 32 338
rect 2080 266 2144 338
rect -32 338 32 482
rect 2080 338 2144 482
rect -32 482 32 554
rect 2080 482 2144 554
<< pdcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 832 68 864 86
rect 832 86 864 104
rect 864 68 928 86
rect 864 86 928 104
rect 928 68 960 86
rect 928 86 960 104
rect 1024 68 1056 86
rect 1024 86 1056 104
rect 1056 68 1120 86
rect 1056 86 1120 104
rect 1120 68 1152 86
rect 1120 86 1152 104
rect 1216 68 1248 86
rect 1216 86 1248 104
rect 1248 68 1312 86
rect 1248 86 1312 104
rect 1312 68 1344 86
rect 1312 86 1344 104
rect 1408 68 1440 86
rect 1408 86 1440 104
rect 1440 68 1504 86
rect 1440 86 1504 104
rect 1504 68 1536 86
rect 1504 86 1536 104
rect 448 284 480 302
rect 448 302 480 320
rect 480 284 544 302
rect 480 302 544 320
rect 544 284 576 302
rect 544 302 576 320
rect 640 284 672 302
rect 640 302 672 320
rect 672 284 736 302
rect 672 302 736 320
rect 736 284 768 302
rect 736 302 768 320
rect 832 284 864 302
rect 832 302 864 320
rect 864 284 928 302
rect 864 302 928 320
rect 928 284 960 302
rect 928 302 960 320
rect 1024 284 1056 302
rect 1024 302 1056 320
rect 1056 284 1120 302
rect 1056 302 1120 320
rect 1120 284 1152 302
rect 1120 302 1152 320
rect 1216 284 1248 302
rect 1216 302 1248 320
rect 1248 284 1312 302
rect 1248 302 1312 320
rect 1312 284 1344 302
rect 1312 302 1344 320
rect 1408 284 1440 302
rect 1408 302 1440 320
rect 1440 284 1504 302
rect 1440 302 1504 320
rect 1504 284 1536 302
rect 1504 302 1536 320
rect 448 500 480 518
rect 448 518 480 536
rect 480 500 544 518
rect 480 518 544 536
rect 544 500 576 518
rect 544 518 576 536
rect 640 500 672 518
rect 640 518 672 536
rect 672 500 736 518
rect 672 518 736 536
rect 736 500 768 518
rect 736 518 768 536
rect 832 500 864 518
rect 832 518 864 536
rect 864 500 928 518
rect 864 518 928 536
rect 928 500 960 518
rect 928 518 960 536
rect 1024 500 1056 518
rect 1024 518 1056 536
rect 1056 500 1120 518
rect 1056 518 1120 536
rect 1120 500 1152 518
rect 1120 518 1152 536
rect 1216 500 1248 518
rect 1216 518 1248 536
rect 1248 500 1312 518
rect 1248 518 1312 536
rect 1312 500 1344 518
rect 1312 518 1344 536
rect 1408 500 1440 518
rect 1408 518 1440 536
rect 1440 500 1504 518
rect 1440 518 1504 536
rect 1504 500 1536 518
rect 1504 518 1536 536
<< nwell >>
rect -184 -124 2296 728
<< labels >>
flabel locali s 1760 338 1824 482 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 1568 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 2016 266 2208 338 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 266 1568 338 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2112 590
<< end >>
