magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1344 459
<< pdiff >>
rect 416 45 800 117
rect 416 117 800 198
rect 416 198 800 270
rect 416 270 800 351
rect 416 351 800 423
<< ntap >>
rect -96 -36 96 45
rect 1248 -36 1440 45
rect -96 45 96 117
rect 1248 45 1440 117
rect -96 117 96 198
rect 1248 117 1440 198
rect -96 198 96 270
rect 1248 198 1440 270
rect -96 270 96 351
rect 1248 270 1440 351
rect -96 351 96 423
rect 1248 351 1440 423
rect -96 423 96 504
rect 1248 423 1440 504
<< poly >>
rect 352 -18 1056 27
rect 352 135 1056 180
rect 352 288 1056 333
rect 352 441 1056 486
rect 992 117 1056 198
rect 992 198 1056 270
rect 992 270 1056 351
<< locali >>
rect 992 270 1056 351
rect -96 -36 96 45
rect 1248 -36 1440 45
rect -96 45 96 117
rect 288 45 800 117
rect 288 45 800 117
rect 1248 45 1440 117
rect -96 117 96 198
rect 288 117 352 198
rect 992 117 1056 198
rect 1248 117 1440 198
rect -96 198 96 270
rect 1248 198 1440 270
rect 288 198 352 270
rect 416 198 800 270
rect 416 198 800 270
rect 992 198 1056 270
rect 1248 198 1440 270
rect -96 270 96 351
rect 288 270 352 351
rect 992 270 1056 351
rect 1248 270 1440 351
rect -96 351 96 423
rect 288 351 800 423
rect 1248 351 1440 423
rect -96 423 96 504
rect 1248 423 1440 504
<< pcontact >>
rect 1002 137 1045 157
rect 1002 157 1045 177
rect 1002 177 1045 197
rect 1002 198 1045 216
rect 1002 216 1045 234
rect 1002 234 1045 252
rect 1002 252 1045 270
rect 1002 270 1045 290
rect 1002 290 1045 310
rect 1002 310 1045 330
<< ntapc >>
rect -32 45 32 117
rect 1312 45 1376 117
rect -32 117 32 198
rect 1312 117 1376 198
rect -32 198 32 270
rect 1312 198 1376 270
rect -32 270 32 351
rect 1312 270 1376 351
rect -32 351 32 423
rect 1312 351 1376 423
<< pdcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 448 216 480 234
rect 448 234 480 252
rect 480 216 544 234
rect 480 234 544 252
rect 544 216 576 234
rect 544 234 576 252
rect 640 216 672 234
rect 640 234 672 252
rect 672 216 736 234
rect 672 234 736 252
rect 736 216 768 234
rect 736 234 768 252
rect 448 369 480 387
rect 448 387 480 405
rect 480 369 544 387
rect 480 387 544 405
rect 544 369 576 387
rect 544 387 576 405
rect 640 369 672 387
rect 640 387 672 405
rect 672 369 736 387
rect 672 387 736 405
rect 736 369 768 387
rect 736 387 768 405
<< nwell >>
rect -184 -124 1528 592
<< labels >>
flabel locali s 992 270 1056 351 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 800 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1248 198 1440 270 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 198 800 270 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1344 459
<< end >>
