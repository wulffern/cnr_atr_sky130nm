magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1152 585
<< pdiff >>
rect 416 45 608 117
rect 416 117 608 261
rect 416 261 608 333
rect 416 333 608 477
rect 416 477 608 549
<< ntap >>
rect -96 -36 96 45
rect 1056 -36 1248 45
rect -96 45 96 117
rect 1056 45 1248 117
rect -96 117 96 261
rect 1056 117 1248 261
rect -96 261 96 333
rect 1056 261 1248 333
rect -96 333 96 477
rect 1056 333 1248 477
rect -96 477 96 549
rect 1056 477 1248 549
rect -96 549 96 630
rect 1056 549 1248 630
<< poly >>
rect 352 -18 864 27
rect 352 135 864 243
rect 352 351 864 459
rect 352 567 864 612
rect 800 117 864 261
rect 800 261 864 333
rect 800 333 864 477
<< locali >>
rect 800 333 864 477
rect -96 -36 96 45
rect 1056 -36 1248 45
rect -96 45 96 117
rect 288 45 608 117
rect 288 45 608 117
rect 1056 45 1248 117
rect -96 117 96 261
rect 288 117 352 261
rect 800 117 864 261
rect 1056 117 1248 261
rect -96 261 96 333
rect 1056 261 1248 333
rect 288 261 352 333
rect 416 261 608 333
rect 416 261 608 333
rect 800 261 864 333
rect 1056 261 1248 333
rect -96 333 96 477
rect 288 333 352 477
rect 800 333 864 477
rect 1056 333 1248 477
rect -96 477 96 549
rect 288 477 608 549
rect 1056 477 1248 549
rect -96 549 96 630
rect 1056 549 1248 630
<< pcontact >>
rect 810 153 853 189
rect 810 189 853 225
rect 810 225 853 261
rect 810 261 853 279
rect 810 279 853 297
rect 810 297 853 315
rect 810 315 853 333
rect 810 333 853 369
rect 810 369 853 405
rect 810 405 853 441
<< ntapc >>
rect -32 45 32 117
rect 1120 45 1184 117
rect -32 117 32 261
rect 1120 117 1184 261
rect -32 261 32 333
rect 1120 261 1184 333
rect -32 333 32 477
rect 1120 333 1184 477
rect -32 477 32 549
rect 1120 477 1184 549
<< pdcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 448 279 480 297
rect 448 297 480 315
rect 480 279 544 297
rect 480 297 544 315
rect 544 279 576 297
rect 544 297 576 315
rect 448 495 480 513
rect 448 513 480 531
rect 480 495 544 513
rect 480 513 544 531
rect 544 495 576 513
rect 544 513 576 531
<< nwell >>
rect -184 -124 1336 718
<< labels >>
flabel locali s 800 333 864 477 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 608 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1056 261 1248 333 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 261 608 333 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 585
<< end >>
