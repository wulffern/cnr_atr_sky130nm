magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 2112 873
<< pdiff >>
rect 416 45 1568 117
rect 416 117 1568 405
rect 416 405 1568 477
rect 416 477 1568 765
rect 416 765 1568 837
<< ntap >>
rect -96 -36 96 45
rect 2016 -36 2208 45
rect -96 45 96 117
rect 2016 45 2208 117
rect -96 117 96 405
rect 2016 117 2208 405
rect -96 405 96 477
rect 2016 405 2208 477
rect -96 477 96 765
rect 2016 477 2208 765
rect -96 765 96 837
rect 2016 765 2208 837
rect -96 837 96 918
rect 2016 837 2208 918
<< poly >>
rect 352 -18 1824 27
rect 352 135 1824 387
rect 352 495 1824 747
rect 352 855 1824 900
rect 1760 117 1824 405
rect 1760 405 1824 477
rect 1760 477 1824 765
<< locali >>
rect 1760 477 1824 765
rect -96 -36 96 45
rect 2016 -36 2208 45
rect -96 45 96 117
rect 288 45 1568 117
rect 288 45 1568 117
rect 2016 45 2208 117
rect -96 117 96 405
rect 288 117 352 405
rect 1760 117 1824 405
rect 2016 117 2208 405
rect -96 405 96 477
rect 2016 405 2208 477
rect 288 405 352 477
rect 416 405 1568 477
rect 416 405 1568 477
rect 1760 405 1824 477
rect 2016 405 2208 477
rect -96 477 96 765
rect 288 477 352 765
rect 1760 477 1824 765
rect 2016 477 2208 765
rect -96 765 96 837
rect 288 765 1568 837
rect 2016 765 2208 837
rect -96 837 96 918
rect 2016 837 2208 918
<< pcontact >>
rect 1770 189 1813 261
rect 1770 261 1813 333
rect 1770 333 1813 405
rect 1770 405 1813 423
rect 1770 423 1813 441
rect 1770 441 1813 459
rect 1770 459 1813 477
rect 1770 477 1813 549
rect 1770 549 1813 621
rect 1770 621 1813 693
<< ntapc >>
rect -32 45 32 117
rect 2080 45 2144 117
rect -32 117 32 405
rect 2080 117 2144 405
rect -32 405 32 477
rect 2080 405 2144 477
rect -32 477 32 765
rect 2080 477 2144 765
rect -32 765 32 837
rect 2080 765 2144 837
<< pdcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 832 63 864 81
rect 832 81 864 99
rect 864 63 928 81
rect 864 81 928 99
rect 928 63 960 81
rect 928 81 960 99
rect 1024 63 1056 81
rect 1024 81 1056 99
rect 1056 63 1120 81
rect 1056 81 1120 99
rect 1120 63 1152 81
rect 1120 81 1152 99
rect 1216 63 1248 81
rect 1216 81 1248 99
rect 1248 63 1312 81
rect 1248 81 1312 99
rect 1312 63 1344 81
rect 1312 81 1344 99
rect 1408 63 1440 81
rect 1408 81 1440 99
rect 1440 63 1504 81
rect 1440 81 1504 99
rect 1504 63 1536 81
rect 1504 81 1536 99
rect 448 423 480 441
rect 448 441 480 459
rect 480 423 544 441
rect 480 441 544 459
rect 544 423 576 441
rect 544 441 576 459
rect 640 423 672 441
rect 640 441 672 459
rect 672 423 736 441
rect 672 441 736 459
rect 736 423 768 441
rect 736 441 768 459
rect 832 423 864 441
rect 832 441 864 459
rect 864 423 928 441
rect 864 441 928 459
rect 928 423 960 441
rect 928 441 960 459
rect 1024 423 1056 441
rect 1024 441 1056 459
rect 1056 423 1120 441
rect 1056 441 1120 459
rect 1120 423 1152 441
rect 1120 441 1152 459
rect 1216 423 1248 441
rect 1216 441 1248 459
rect 1248 423 1312 441
rect 1248 441 1312 459
rect 1312 423 1344 441
rect 1312 441 1344 459
rect 1408 423 1440 441
rect 1408 441 1440 459
rect 1440 423 1504 441
rect 1440 441 1504 459
rect 1504 423 1536 441
rect 1504 441 1536 459
rect 448 783 480 801
rect 448 801 480 819
rect 480 783 544 801
rect 480 801 544 819
rect 544 783 576 801
rect 544 801 576 819
rect 640 783 672 801
rect 640 801 672 819
rect 672 783 736 801
rect 672 801 736 819
rect 736 783 768 801
rect 736 801 768 819
rect 832 783 864 801
rect 832 801 864 819
rect 864 783 928 801
rect 864 801 928 819
rect 928 783 960 801
rect 928 801 960 819
rect 1024 783 1056 801
rect 1024 801 1056 819
rect 1056 783 1120 801
rect 1056 801 1120 819
rect 1120 783 1152 801
rect 1120 801 1152 819
rect 1216 783 1248 801
rect 1216 801 1248 819
rect 1248 783 1312 801
rect 1248 801 1312 819
rect 1312 783 1344 801
rect 1312 801 1344 819
rect 1408 783 1440 801
rect 1408 801 1440 819
rect 1440 783 1504 801
rect 1440 801 1504 819
rect 1504 783 1536 801
rect 1504 801 1536 819
<< nwell >>
rect -184 -124 2296 1006
<< labels >>
flabel locali s 1760 477 1824 765 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 1568 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 2016 405 2208 477 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 405 1568 477 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2112 873
<< end >>
