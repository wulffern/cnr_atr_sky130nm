magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1728 2025
<< ndiff >>
rect 416 45 1184 117
rect 416 117 1184 981
rect 416 981 1184 1053
rect 416 1053 1184 1917
rect 416 1917 1184 1989
<< ptap >>
rect -96 -36 96 45
rect 1632 -36 1824 45
rect -96 45 96 117
rect 1632 45 1824 117
rect -96 117 96 981
rect 1632 117 1824 981
rect -96 981 96 1053
rect 1632 981 1824 1053
rect -96 1053 96 1917
rect 1632 1053 1824 1917
rect -96 1917 96 1989
rect 1632 1917 1824 1989
rect -96 1989 96 2070
rect 1632 1989 1824 2070
<< poly >>
rect 352 -18 1440 27
rect 352 135 1440 963
rect 352 1071 1440 1899
rect 352 2007 1440 2052
rect 1376 117 1440 981
rect 1376 981 1440 1053
rect 1376 1053 1440 1917
<< locali >>
rect 1376 1053 1440 1917
rect -96 -36 96 45
rect 1632 -36 1824 45
rect -96 45 96 117
rect 288 45 1184 117
rect 288 45 1184 117
rect 1632 45 1824 117
rect -96 117 96 981
rect 288 117 352 981
rect 1376 117 1440 981
rect 1632 117 1824 981
rect -96 981 96 1053
rect 1632 981 1824 1053
rect 288 981 352 1053
rect 416 981 1184 1053
rect 416 981 1184 1053
rect 1376 981 1440 1053
rect 1632 981 1824 1053
rect -96 1053 96 1917
rect 288 1053 352 1917
rect 1376 1053 1440 1917
rect 1632 1053 1824 1917
rect -96 1917 96 1989
rect 288 1917 1184 1989
rect 1632 1917 1824 1989
rect -96 1989 96 2070
rect 1632 1989 1824 2070
<< pcontact >>
rect 1386 333 1429 549
rect 1386 549 1429 765
rect 1386 765 1429 981
rect 1386 981 1429 999
rect 1386 999 1429 1017
rect 1386 1017 1429 1035
rect 1386 1035 1429 1053
rect 1386 1053 1429 1269
rect 1386 1269 1429 1485
rect 1386 1485 1429 1701
<< ptapc >>
rect -32 45 32 117
rect 1696 45 1760 117
rect -32 117 32 981
rect 1696 117 1760 981
rect -32 981 32 1053
rect 1696 981 1760 1053
rect -32 1053 32 1917
rect 1696 1053 1760 1917
rect -32 1917 32 1989
rect 1696 1917 1760 1989
<< ndcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 832 63 864 81
rect 832 81 864 99
rect 864 63 928 81
rect 864 81 928 99
rect 928 63 960 81
rect 928 81 960 99
rect 1024 63 1056 81
rect 1024 81 1056 99
rect 1056 63 1120 81
rect 1056 81 1120 99
rect 1120 63 1152 81
rect 1120 81 1152 99
rect 448 999 480 1017
rect 448 1017 480 1035
rect 480 999 544 1017
rect 480 1017 544 1035
rect 544 999 576 1017
rect 544 1017 576 1035
rect 640 999 672 1017
rect 640 1017 672 1035
rect 672 999 736 1017
rect 672 1017 736 1035
rect 736 999 768 1017
rect 736 1017 768 1035
rect 832 999 864 1017
rect 832 1017 864 1035
rect 864 999 928 1017
rect 864 1017 928 1035
rect 928 999 960 1017
rect 928 1017 960 1035
rect 1024 999 1056 1017
rect 1024 1017 1056 1035
rect 1056 999 1120 1017
rect 1056 1017 1120 1035
rect 1120 999 1152 1017
rect 1120 1017 1152 1035
rect 448 1935 480 1953
rect 448 1953 480 1971
rect 480 1935 544 1953
rect 480 1953 544 1971
rect 544 1935 576 1953
rect 544 1953 576 1971
rect 640 1935 672 1953
rect 640 1953 672 1971
rect 672 1935 736 1953
rect 672 1953 736 1971
rect 736 1935 768 1953
rect 736 1953 768 1971
rect 832 1935 864 1953
rect 832 1953 864 1971
rect 864 1935 928 1953
rect 864 1953 928 1971
rect 928 1935 960 1953
rect 928 1953 960 1971
rect 1024 1935 1056 1953
rect 1024 1953 1056 1971
rect 1056 1935 1120 1953
rect 1056 1953 1120 1971
rect 1120 1935 1152 1953
rect 1120 1953 1152 1971
<< pwell >>
rect -184 -124 1912 2158
<< labels >>
flabel locali s 1376 1053 1440 1917 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 1184 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1632 981 1824 1053 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 981 1184 1053 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1728 2025
<< end >>
