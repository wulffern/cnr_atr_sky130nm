magic
tech sky130B
magscale 1 2
timestamp 1712008800
<< checkpaint >>
rect 0 0 1728 459
<< ndiff >>
rect 416 45 1184 117
rect 416 117 1184 198
rect 416 198 1184 270
rect 416 270 1184 351
rect 416 351 1184 423
<< ptap >>
rect -96 -36 96 45
rect 1632 -36 1824 45
rect -96 45 96 117
rect 1632 45 1824 117
rect -96 117 96 198
rect 1632 117 1824 198
rect -96 198 96 270
rect 1632 198 1824 270
rect -96 270 96 351
rect 1632 270 1824 351
rect -96 351 96 423
rect 1632 351 1824 423
rect -96 423 96 504
rect 1632 423 1824 504
<< poly >>
rect 352 -18 1440 27
rect 352 135 1440 180
rect 352 288 1440 333
rect 352 441 1440 486
rect 1376 117 1440 198
rect 1376 198 1440 270
rect 1376 270 1440 351
<< locali >>
rect 1376 270 1440 351
rect -96 -36 96 45
rect 1632 -36 1824 45
rect -96 45 96 117
rect 288 45 1184 117
rect 288 45 1184 117
rect 1632 45 1824 117
rect -96 117 96 198
rect 288 117 352 198
rect 1376 117 1440 198
rect 1632 117 1824 198
rect -96 198 96 270
rect 1632 198 1824 270
rect 288 198 352 270
rect 416 198 1184 270
rect 416 198 1184 270
rect 1376 198 1440 270
rect 1632 198 1824 270
rect -96 270 96 351
rect 288 270 352 351
rect 1376 270 1440 351
rect 1632 270 1824 351
rect -96 351 96 423
rect 288 351 1184 423
rect 1632 351 1824 423
rect -96 423 96 504
rect 1632 423 1824 504
<< pcontact >>
rect 1386 137 1429 157
rect 1386 157 1429 177
rect 1386 177 1429 197
rect 1386 198 1429 216
rect 1386 216 1429 234
rect 1386 234 1429 252
rect 1386 252 1429 270
rect 1386 270 1429 290
rect 1386 290 1429 310
rect 1386 310 1429 330
<< ptapc >>
rect -32 45 32 117
rect 1696 45 1760 117
rect -32 117 32 198
rect 1696 117 1760 198
rect -32 198 32 270
rect 1696 198 1760 270
rect -32 270 32 351
rect 1696 270 1760 351
rect -32 351 32 423
rect 1696 351 1760 423
<< ndcontact >>
rect 448 63 480 81
rect 448 81 480 99
rect 480 63 544 81
rect 480 81 544 99
rect 544 63 576 81
rect 544 81 576 99
rect 640 63 672 81
rect 640 81 672 99
rect 672 63 736 81
rect 672 81 736 99
rect 736 63 768 81
rect 736 81 768 99
rect 832 63 864 81
rect 832 81 864 99
rect 864 63 928 81
rect 864 81 928 99
rect 928 63 960 81
rect 928 81 960 99
rect 1024 63 1056 81
rect 1024 81 1056 99
rect 1056 63 1120 81
rect 1056 81 1120 99
rect 1120 63 1152 81
rect 1120 81 1152 99
rect 448 216 480 234
rect 448 234 480 252
rect 480 216 544 234
rect 480 234 544 252
rect 544 216 576 234
rect 544 234 576 252
rect 640 216 672 234
rect 640 234 672 252
rect 672 216 736 234
rect 672 234 736 252
rect 736 216 768 234
rect 736 234 768 252
rect 832 216 864 234
rect 832 234 864 252
rect 864 216 928 234
rect 864 234 928 252
rect 928 216 960 234
rect 928 234 960 252
rect 1024 216 1056 234
rect 1024 234 1056 252
rect 1056 216 1120 234
rect 1056 234 1120 252
rect 1120 216 1152 234
rect 1120 234 1152 252
rect 448 369 480 387
rect 448 387 480 405
rect 480 369 544 387
rect 480 387 544 405
rect 544 369 576 387
rect 544 387 576 405
rect 640 369 672 387
rect 640 387 672 405
rect 672 369 736 387
rect 672 387 736 405
rect 736 369 768 387
rect 736 387 768 405
rect 832 369 864 387
rect 832 387 864 405
rect 864 369 928 387
rect 864 387 928 405
rect 928 369 960 387
rect 928 387 960 405
rect 1024 369 1056 387
rect 1024 387 1056 405
rect 1056 369 1120 387
rect 1056 387 1120 405
rect 1120 369 1152 387
rect 1120 387 1152 405
<< pwell >>
rect -184 -124 1912 592
<< labels >>
flabel locali s 1376 270 1440 351 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 45 1184 117 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1632 198 1824 270 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 198 1184 270 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1728 459
<< end >>
