magic
tech sky130B
magscale 1 2
timestamp 1695852000
<< checkpaint >>
rect 0 0 1728 1454
<< ndiff >>
rect 416 50 1184 122
rect 416 122 1184 698
rect 416 698 1184 770
rect 416 770 1184 1346
rect 416 1346 1184 1418
<< ptap >>
rect -96 -36 96 50
rect 1632 -36 1824 50
rect -96 50 96 122
rect 1632 50 1824 122
rect -96 122 96 698
rect 1632 122 1824 698
rect -96 698 96 770
rect 1632 698 1824 770
rect -96 770 96 1346
rect 1632 770 1824 1346
rect -96 1346 96 1418
rect 1632 1346 1824 1418
rect -96 1418 96 1504
rect 1632 1418 1824 1504
<< poly >>
rect 352 -18 1440 32
rect 352 140 1440 680
rect 352 788 1440 1328
rect 352 1436 1440 1486
rect 1376 122 1440 698
rect 1376 698 1440 770
rect 1376 770 1440 1346
<< locali >>
rect 1376 770 1440 1346
rect -96 -36 96 50
rect 1632 -36 1824 50
rect -96 50 96 122
rect 288 50 1184 122
rect 288 50 1184 122
rect 1632 50 1824 122
rect -96 122 96 698
rect 288 122 352 698
rect 1376 122 1440 698
rect 1632 122 1824 698
rect -96 698 96 770
rect 1632 698 1824 770
rect 288 698 352 770
rect 416 698 1184 770
rect 416 698 1184 770
rect 1376 698 1440 770
rect 1632 698 1824 770
rect -96 770 96 1346
rect 288 770 352 1346
rect 1376 770 1440 1346
rect 1632 770 1824 1346
rect -96 1346 96 1418
rect 288 1346 1184 1418
rect 1632 1346 1824 1418
rect -96 1418 96 1504
rect 1632 1418 1824 1504
<< pcontact >>
rect 1386 266 1429 410
rect 1386 410 1429 554
rect 1386 554 1429 698
rect 1386 698 1429 716
rect 1386 716 1429 734
rect 1386 734 1429 752
rect 1386 752 1429 770
rect 1386 770 1429 914
rect 1386 914 1429 1058
rect 1386 1058 1429 1202
<< ptapc >>
rect -32 50 32 122
rect 1696 50 1760 122
rect -32 122 32 698
rect 1696 122 1760 698
rect -32 698 32 770
rect 1696 698 1760 770
rect -32 770 32 1346
rect 1696 770 1760 1346
rect -32 1346 32 1418
rect 1696 1346 1760 1418
<< ndcontact >>
rect 448 68 480 86
rect 448 86 480 104
rect 480 68 544 86
rect 480 86 544 104
rect 544 68 576 86
rect 544 86 576 104
rect 640 68 672 86
rect 640 86 672 104
rect 672 68 736 86
rect 672 86 736 104
rect 736 68 768 86
rect 736 86 768 104
rect 832 68 864 86
rect 832 86 864 104
rect 864 68 928 86
rect 864 86 928 104
rect 928 68 960 86
rect 928 86 960 104
rect 1024 68 1056 86
rect 1024 86 1056 104
rect 1056 68 1120 86
rect 1056 86 1120 104
rect 1120 68 1152 86
rect 1120 86 1152 104
rect 448 716 480 734
rect 448 734 480 752
rect 480 716 544 734
rect 480 734 544 752
rect 544 716 576 734
rect 544 734 576 752
rect 640 716 672 734
rect 640 734 672 752
rect 672 716 736 734
rect 672 734 736 752
rect 736 716 768 734
rect 736 734 768 752
rect 832 716 864 734
rect 832 734 864 752
rect 864 716 928 734
rect 864 734 928 752
rect 928 716 960 734
rect 928 734 960 752
rect 1024 716 1056 734
rect 1024 734 1056 752
rect 1056 716 1120 734
rect 1056 734 1120 752
rect 1120 716 1152 734
rect 1120 734 1152 752
rect 448 1364 480 1382
rect 448 1382 480 1400
rect 480 1364 544 1382
rect 480 1382 544 1400
rect 544 1364 576 1382
rect 544 1382 576 1400
rect 640 1364 672 1382
rect 640 1382 672 1400
rect 672 1364 736 1382
rect 672 1382 736 1400
rect 736 1364 768 1382
rect 736 1382 768 1400
rect 832 1364 864 1382
rect 832 1382 864 1400
rect 864 1364 928 1382
rect 864 1382 928 1400
rect 928 1364 960 1382
rect 928 1382 960 1400
rect 1024 1364 1056 1382
rect 1024 1382 1056 1400
rect 1056 1364 1120 1382
rect 1056 1382 1120 1400
rect 1120 1364 1152 1382
rect 1120 1382 1152 1400
<< pwell >>
rect -184 -124 1912 1592
<< labels >>
flabel locali s 1376 770 1440 1346 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 288 50 1184 122 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 1632 698 1824 770 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 416 698 1184 770 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1728 1454
<< end >>
