
//-------------------------------------------------------------
// CNRATR_PCH_2C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_2C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_2C2F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_2C2F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_2C4F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_2C4F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_2C8F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_2C8F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_2C12F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_2C12F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_4C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_4C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_4C2F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_4C2F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_4C4F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_4C4F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_4C8F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_4C8F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_4C12F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_4C12F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_8C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_8C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_8C2F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_8C2F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_8C4F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_8C4F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_8C8F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_8C8F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_8C12F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_8C12F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_12C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_12C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_12C2F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_12C2F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_12C4F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_12C4F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_12C8F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_12C8F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_PCH_12C12F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_PCH_12C12F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_2C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_2C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_2C2F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_2C2F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_2C4F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_2C4F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_2C8F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_2C8F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_2C12F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_2C12F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_4C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_4C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_4C2F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_4C2F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_4C4F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_4C4F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_4C8F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_4C8F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_4C12F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_4C12F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_8C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_8C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_8C2F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_8C2F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_8C4F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_8C4F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_8C8F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_8C8F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_8C12F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_8C12F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_12C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_12C1F2(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_12C2F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_12C2F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_12C4F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_12C4F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_12C8F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_12C8F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule

//-------------------------------------------------------------
// CNRATR_NCH_12C12F0 <class 'cicpy.core.layoutcell.LayoutCell'>
//-------------------------------------------------------------
module CNRATR_NCH_12C12F0(D,G,S,B);
input logic G;
input logic S;
input logic B;
input logic D;
endmodule
